module z_sign_extend_17_32(in, out);
	input [16:0] in;
	output [31:0] out;
	
	assign out[16:0] = in;
	genvar i;
	generate
		for (i=17; i<32; i=i+1) begin: loop1
			assign out[i] = in[16];
		end
	endgenerate
endmodule