module multdiv(data_operandA, data_operandB, ctrl_MULT, ctrl_DIV, clock, data_result, data_exception, data_resultRDY);
   input [31:0] data_operandA, data_operandB;
   input ctrl_MULT, ctrl_DIV, clock;
	
   output [31:0] data_result; 
	output data_exception, data_resultRDY;
	
	// opcode (mult/div) memory
	wire writeOpHolder, currentOp;
	or(writeOpHolder, ctrl_MULT, ctrl_DIV);
	reg_1 opHolder(ctrl_MULT, clock, 1'b1, writeOpHolder, currentOp);
	
	wire [31:0] hold_dataA_mult, hold_dataB_mult;
	
	reg_32 storeA(data_operandA, clock, 1'b1, ctrl_MULT, hold_dataA_mult);
	reg_32 storeB(data_operandB, clock, 1'b1, ctrl_MULT, hold_dataB_mult);
	
	
	// mult
	wire [2:0] counter_wire_mult;
   wire [31:0] mult_data_result;
	wire mult_data_exception;
	counter_reg3 counter_mult(clock, writeOpHolder, 1'b1, counter_wire_mult);
	wallace w1(mult_data_result, hold_dataA_mult, hold_dataB_mult, ctrl_MULT, mult_data_exception);
	
	
	// Create registers to store data_operandA and data_operandB

	
	
	// div
	
	wire [33:0] counter_wire_div;
	wire [32:0] pre_div_data_result;
	wire [31:0] pos_div_data_result, neg_div_data_result, div_data_result;
	wire div_data_exception;
	wire [31:0] pos_data_operandA, pos_data_operandB;
	counter_reg34 counter_div(clock, writeOpHolder, 1'b1, counter_wire_div);
	abs32 abs1(pos_data_operandA, data_operandA);
	abs32 abs2(pos_data_operandB, data_operandB);
	
	wire [31:0] hold_pos_data_operandA_div, hold_pos_data_operandB_div;	
	reg_32 storeAdiv(pos_data_operandA, clock, 1'b1, ctrl_DIV, hold_pos_data_operandA_div);
	reg_32 storeBdiv(pos_data_operandB, clock, 1'b1, ctrl_DIV, hold_pos_data_operandB_div);
	
	divider d1(hold_pos_data_operandA_div, hold_pos_data_operandB_div, counter_wire_div, ctrl_DIV, clock, 1'b1, pre_div_data_result, div_data_exception);
	
	// post divider logic
	assign pos_div_data_result = pre_div_data_result[32:1];
	wire keepResult;
	isNegRes ng1(keepResult, data_operandA[31], data_operandB[31]);
	twoscomp32 negativeRes(neg_div_data_result, pos_div_data_result);
	assign div_data_result = keepResult ? pos_div_data_result : neg_div_data_result;
	
	
	
	// MUX AT THE END
	//assign data_exception
	assign data_result = currentOp ? mult_data_result : div_data_result;
	assign data_exception = currentOp ? mult_data_exception : div_data_exception;
	assign data_resultRDY = currentOp ? counter_wire_mult[2] : counter_wire_div[33];
	
	//	// Your code here
	//	wire [2:0] counter_wire_mult;
	//	counter_reg3 counter_mult(clock, ctrl_MULT, 1'b1, counter_wire_mult);
	//	wallace m1(data_result, pos_data_operandA, pos_data_operandB, ctrl_MULT, data_exception);
	//	
endmodule

module divider(dividend, divisor, counterWire, l_stg, clk, enable, data_result, de);
    // Initialize inputs, both dividend and divisor MUST BE positive
    input [31:0] dividend, divisor;
	 input [33:0] counterWire;
    input l_stg, clk, enable;

    // Initialize outputs
    output [32:0] data_result;
    output de;

    // Initialize wires
    wire [63:0] curr_regval, post_subtract, post_shift, next_regval;
    wire [31:0] sub_res, most_sigbits, added_1, least_sigbits;
    wire perform_subtract;
    
    // Subtract divisor from top half. 
    wire cout_sub;
    cselect_adder_32 subtract_op(curr_regval[63:32], ~divisor, 1'b1, cout_sub, sub_res);
	 // if the result from LHS-divisor is negative, we must NOT subtract
    assign perform_subtract = sub_res[31];

    assign most_sigbits = perform_subtract ? curr_regval[63:32] : sub_res;
    
	 // Added_1 represents the rhs where u add 1 if u are able to successfully subtract
    assign added_1[31:1] = curr_regval[31:1];
    assign added_1[0] = 1'b1;

    // Mux between subtract divisor or not subtract divisor.
    assign least_sigbits = perform_subtract ? curr_regval[31:0] : added_1; 

    // After subtract/no subtract
    assign post_subtract[63:32] = most_sigbits;
    assign post_subtract[31:0] = least_sigbits;

    // Left Shift.
	 
	 assign post_shift = post_subtract << 1;
	 
	 wire [63:0] post_shift_final;
	 assign post_shift_final = counterWire[33] ? post_subtract : post_shift;

    assign next_regval[63:32] = l_stg ? 32'b0 : post_shift_final[63:32];
    assign next_regval[31:0] = l_stg ? dividend : post_shift_final[31:0];
	 
	 // if counter register equals 1 then just subtract if possible without shifting
	 //wire cout_sub_two;
	 //wire [31:0] sub_res_two;
	 //cselect_adder_32 subtract_two(next_regval[63:32], ~divisor, 1'b1, cout_sub_two, sub_res_two);
	 //assign perform_subtract_two = sub_res_two[31];

    reg_64 quiotient(next_regval, clk, 1'b1, enable, curr_regval);

    assign data_result = curr_regval[32:0];
    //assign de = divisor ? 1'b0 :1'b1;
	 assign de = 1'b0;
endmodule

// Counter Registers 
module counter_reg(clk, reset, enable, out);
	input reset, clk, enable;
	
	wire [32:0] reg_curr_val, reg_next_val, shifted_val, register_value;
	output [32:0] out;
	
	// Shift register value in count step
   l_shift_1 y1(register_value, shifted_val);

	assign out = reg_curr_val;
	assign reg_next_val = reset ? 33'b1 : shifted_val;
	
	reg_32 reg0_31(reg_next_val[31:0], clk, 1'b1, enable, reg_curr_val[31:0]);
	reg_1 reg32(reg_next_val[32], clk, 1'b1, enable, reg_curr_val[32]);
endmodule

module counter_reg3(clk, reset, enable, out);
	input reset, clk, enable;
	
	wire [2:0] reg_curr_val, reg_next_val, shifted_val;
	output [2:0] out;
	
	// Shift register value in count step
   l_shift_1 r(reg_curr_val, shifted_val);

	assign out = reg_curr_val;
	assign reg_next_val = reset ? 3'b001 : shifted_val;
	
	reg_3 reg3(reg_next_val, clk, 1'b1, enable, reg_curr_val);
endmodule

module counter_reg33(clk, reset, enable, out);
	input reset, clk, enable;
	
	wire [32:0] reg_curr_val, reg_next_val, shifted_val;
	output [32:0] out;
	
	// Shift register value in count step
	assign shifted_val = reg_curr_val << 1;

	assign out = reg_curr_val;
	assign reg_next_val = reset ? 33'b000000000000000000000000000000001 : shifted_val;
	
	reg_33 reg33(reg_next_val, clk, 1'b1, enable, reg_curr_val);
endmodule

module counter_reg34(clk, reset, enable, out);
	input reset, clk, enable;
	
	wire [33:0] reg_curr_val, reg_next_val, shifted_val;
	output [33:0] out;
	
	// Shift register value in count step
	assign shifted_val = reg_curr_val << 1;

	assign out = reg_curr_val;
	assign reg_next_val = reset ? 34'b0000000000000000000000000000000001 : shifted_val;
	
	reg_34 reg34(reg_next_val, clk, 1'b1, enable, reg_curr_val);
endmodule

module isNegRes(out, a, b);
	input a, b;
	output out;
	
	wire out1, out2;

	and and1(out1, a, b);
	and and2(out2,~a, ~b);
	
	or(out,out1,out2);
endmodule

module full_adder_md(s, cout, in1, in2, cin);
	input in1, in2, cin;
	output cout, s;
	
	wire out_xor1, out_and1, out_and2;
	
	
	xor xor1(out_xor1, in1, in2);
	and and1(out_and1, in1, in2);
	xor xor2(s, out_xor1, cin);
	and and2(out_and2, out_xor1, cin);
	or or1(cout, out_and1, out_and2);
endmodule

module wallace (data_result, data_operandA, data_operandB, ctrl_MULT, data_exception);

	input [31:0] data_operandA, data_operandB;
	input ctrl_MULT;

	output [31:0] data_result;
	output data_exception;

	// TODO
	assign data_exception = 1'b0;

	wire w_stg_0_0_0, w_stg_0_0_1, w_stg_0_0_2, w_stg_0_0_3, w_stg_0_0_4, w_stg_0_0_5, w_stg_0_0_6, w_stg_0_0_7, w_stg_0_0_8, w_stg_0_0_9, w_stg_0_0_10, w_stg_0_0_11, w_stg_0_0_12, w_stg_0_0_13, w_stg_0_0_14, w_stg_0_0_15, w_stg_0_0_16, w_stg_0_0_17, w_stg_0_0_18, w_stg_0_0_19, w_stg_0_0_20, w_stg_0_0_21, w_stg_0_0_22, w_stg_0_0_23, w_stg_0_0_24, w_stg_0_0_25, w_stg_0_0_26, w_stg_0_0_27, w_stg_0_0_28, w_stg_0_0_29, w_stg_0_0_30, w_stg_0_0_31, w_stg_0_1_1, w_stg_0_1_2, w_stg_0_1_3, w_stg_0_1_4, w_stg_0_1_5, w_stg_0_1_6, w_stg_0_1_7, w_stg_0_1_8, w_stg_0_1_9, w_stg_0_1_10, w_stg_0_1_11, w_stg_0_1_12, w_stg_0_1_13, w_stg_0_1_14, w_stg_0_1_15, w_stg_0_1_16, w_stg_0_1_17, w_stg_0_1_18, w_stg_0_1_19, w_stg_0_1_20, w_stg_0_1_21, w_stg_0_1_22, w_stg_0_1_23, w_stg_0_1_24, w_stg_0_1_25, w_stg_0_1_26, w_stg_0_1_27, w_stg_0_1_28, w_stg_0_1_29, w_stg_0_1_30, w_stg_0_1_31, w_stg_0_1_32, w_stg_0_2_2, w_stg_0_2_3, w_stg_0_2_4, w_stg_0_2_5, w_stg_0_2_6, w_stg_0_2_7, w_stg_0_2_8, w_stg_0_2_9, w_stg_0_2_10, w_stg_0_2_11, w_stg_0_2_12, w_stg_0_2_13, w_stg_0_2_14, w_stg_0_2_15, w_stg_0_2_16, w_stg_0_2_17, w_stg_0_2_18, w_stg_0_2_19, w_stg_0_2_20, w_stg_0_2_21, w_stg_0_2_22, w_stg_0_2_23, w_stg_0_2_24, w_stg_0_2_25, w_stg_0_2_26, w_stg_0_2_27, w_stg_0_2_28, w_stg_0_2_29, w_stg_0_2_30, w_stg_0_2_31, w_stg_0_2_32, w_stg_0_2_33, w_stg_0_3_3, w_stg_0_3_4, w_stg_0_3_5, w_stg_0_3_6, w_stg_0_3_7, w_stg_0_3_8, w_stg_0_3_9, w_stg_0_3_10, w_stg_0_3_11, w_stg_0_3_12, w_stg_0_3_13, w_stg_0_3_14, w_stg_0_3_15, w_stg_0_3_16, w_stg_0_3_17, w_stg_0_3_18, w_stg_0_3_19, w_stg_0_3_20, w_stg_0_3_21, w_stg_0_3_22, w_stg_0_3_23, w_stg_0_3_24, w_stg_0_3_25, w_stg_0_3_26, w_stg_0_3_27, w_stg_0_3_28, w_stg_0_3_29, w_stg_0_3_30, w_stg_0_3_31, w_stg_0_3_32, w_stg_0_3_33, w_stg_0_3_34, w_stg_0_4_4, w_stg_0_4_5, w_stg_0_4_6, w_stg_0_4_7, w_stg_0_4_8, w_stg_0_4_9, w_stg_0_4_10, w_stg_0_4_11, w_stg_0_4_12, w_stg_0_4_13, w_stg_0_4_14, w_stg_0_4_15, w_stg_0_4_16, w_stg_0_4_17, w_stg_0_4_18, w_stg_0_4_19, w_stg_0_4_20, w_stg_0_4_21, w_stg_0_4_22, w_stg_0_4_23, w_stg_0_4_24, w_stg_0_4_25, w_stg_0_4_26, w_stg_0_4_27, w_stg_0_4_28, w_stg_0_4_29, w_stg_0_4_30, w_stg_0_4_31, w_stg_0_4_32, w_stg_0_4_33, w_stg_0_4_34, w_stg_0_4_35, w_stg_0_5_5, w_stg_0_5_6, w_stg_0_5_7, w_stg_0_5_8, w_stg_0_5_9, w_stg_0_5_10, w_stg_0_5_11, w_stg_0_5_12, w_stg_0_5_13, w_stg_0_5_14, w_stg_0_5_15, w_stg_0_5_16, w_stg_0_5_17, w_stg_0_5_18, w_stg_0_5_19, w_stg_0_5_20, w_stg_0_5_21, w_stg_0_5_22, w_stg_0_5_23, w_stg_0_5_24, w_stg_0_5_25, w_stg_0_5_26, w_stg_0_5_27, w_stg_0_5_28, w_stg_0_5_29, w_stg_0_5_30, w_stg_0_5_31, w_stg_0_5_32, w_stg_0_5_33, w_stg_0_5_34, w_stg_0_5_35, w_stg_0_5_36, w_stg_0_6_6, w_stg_0_6_7, w_stg_0_6_8, w_stg_0_6_9, w_stg_0_6_10, w_stg_0_6_11, w_stg_0_6_12, w_stg_0_6_13, w_stg_0_6_14, w_stg_0_6_15, w_stg_0_6_16, w_stg_0_6_17, w_stg_0_6_18, w_stg_0_6_19, w_stg_0_6_20, w_stg_0_6_21, w_stg_0_6_22, w_stg_0_6_23, w_stg_0_6_24, w_stg_0_6_25, w_stg_0_6_26, w_stg_0_6_27, w_stg_0_6_28, w_stg_0_6_29, w_stg_0_6_30, w_stg_0_6_31, w_stg_0_6_32, w_stg_0_6_33, w_stg_0_6_34, w_stg_0_6_35, w_stg_0_6_36, w_stg_0_6_37, w_stg_0_7_7, w_stg_0_7_8, w_stg_0_7_9, w_stg_0_7_10, w_stg_0_7_11, w_stg_0_7_12, w_stg_0_7_13, w_stg_0_7_14, w_stg_0_7_15, w_stg_0_7_16, w_stg_0_7_17, w_stg_0_7_18, w_stg_0_7_19, w_stg_0_7_20, w_stg_0_7_21, w_stg_0_7_22, w_stg_0_7_23, w_stg_0_7_24, w_stg_0_7_25, w_stg_0_7_26, w_stg_0_7_27, w_stg_0_7_28, w_stg_0_7_29, w_stg_0_7_30, w_stg_0_7_31, w_stg_0_7_32, w_stg_0_7_33, w_stg_0_7_34, w_stg_0_7_35, w_stg_0_7_36, w_stg_0_7_37, w_stg_0_7_38, w_stg_0_8_8, w_stg_0_8_9, w_stg_0_8_10, w_stg_0_8_11, w_stg_0_8_12, w_stg_0_8_13, w_stg_0_8_14, w_stg_0_8_15, w_stg_0_8_16, w_stg_0_8_17, w_stg_0_8_18, w_stg_0_8_19, w_stg_0_8_20, w_stg_0_8_21, w_stg_0_8_22, w_stg_0_8_23, w_stg_0_8_24, w_stg_0_8_25, w_stg_0_8_26, w_stg_0_8_27, w_stg_0_8_28, w_stg_0_8_29, w_stg_0_8_30, w_stg_0_8_31, w_stg_0_8_32, w_stg_0_8_33, w_stg_0_8_34, w_stg_0_8_35, w_stg_0_8_36, w_stg_0_8_37, w_stg_0_8_38, w_stg_0_8_39, w_stg_0_9_9, w_stg_0_9_10, w_stg_0_9_11, w_stg_0_9_12, w_stg_0_9_13, w_stg_0_9_14, w_stg_0_9_15, w_stg_0_9_16, w_stg_0_9_17, w_stg_0_9_18, w_stg_0_9_19, w_stg_0_9_20, w_stg_0_9_21, w_stg_0_9_22, w_stg_0_9_23, w_stg_0_9_24, w_stg_0_9_25, w_stg_0_9_26, w_stg_0_9_27, w_stg_0_9_28, w_stg_0_9_29, w_stg_0_9_30, w_stg_0_9_31, w_stg_0_9_32, w_stg_0_9_33, w_stg_0_9_34, w_stg_0_9_35, w_stg_0_9_36, w_stg_0_9_37, w_stg_0_9_38, w_stg_0_9_39, w_stg_0_9_40, w_stg_0_10_10, w_stg_0_10_11, w_stg_0_10_12, w_stg_0_10_13, w_stg_0_10_14, w_stg_0_10_15, w_stg_0_10_16, w_stg_0_10_17, w_stg_0_10_18, w_stg_0_10_19, w_stg_0_10_20, w_stg_0_10_21, w_stg_0_10_22, w_stg_0_10_23, w_stg_0_10_24, w_stg_0_10_25, w_stg_0_10_26, w_stg_0_10_27, w_stg_0_10_28, w_stg_0_10_29, w_stg_0_10_30, w_stg_0_10_31, w_stg_0_10_32, w_stg_0_10_33, w_stg_0_10_34, w_stg_0_10_35, w_stg_0_10_36, w_stg_0_10_37, w_stg_0_10_38, w_stg_0_10_39, w_stg_0_10_40, w_stg_0_10_41, w_stg_0_11_11, w_stg_0_11_12, w_stg_0_11_13, w_stg_0_11_14, w_stg_0_11_15, w_stg_0_11_16, w_stg_0_11_17, w_stg_0_11_18, w_stg_0_11_19, w_stg_0_11_20, w_stg_0_11_21, w_stg_0_11_22, w_stg_0_11_23, w_stg_0_11_24, w_stg_0_11_25, w_stg_0_11_26, w_stg_0_11_27, w_stg_0_11_28, w_stg_0_11_29, w_stg_0_11_30, w_stg_0_11_31, w_stg_0_11_32, w_stg_0_11_33, w_stg_0_11_34, w_stg_0_11_35, w_stg_0_11_36, w_stg_0_11_37, w_stg_0_11_38, w_stg_0_11_39, w_stg_0_11_40, w_stg_0_11_41, w_stg_0_11_42, w_stg_0_12_12, w_stg_0_12_13, w_stg_0_12_14, w_stg_0_12_15, w_stg_0_12_16, w_stg_0_12_17, w_stg_0_12_18, w_stg_0_12_19, w_stg_0_12_20, w_stg_0_12_21, w_stg_0_12_22, w_stg_0_12_23, w_stg_0_12_24, w_stg_0_12_25, w_stg_0_12_26, w_stg_0_12_27, w_stg_0_12_28, w_stg_0_12_29, w_stg_0_12_30, w_stg_0_12_31, w_stg_0_12_32, w_stg_0_12_33, w_stg_0_12_34, w_stg_0_12_35, w_stg_0_12_36, w_stg_0_12_37, w_stg_0_12_38, w_stg_0_12_39, w_stg_0_12_40, w_stg_0_12_41, w_stg_0_12_42, w_stg_0_12_43, w_stg_0_13_13, w_stg_0_13_14, w_stg_0_13_15, w_stg_0_13_16, w_stg_0_13_17, w_stg_0_13_18, w_stg_0_13_19, w_stg_0_13_20, w_stg_0_13_21, w_stg_0_13_22, w_stg_0_13_23, w_stg_0_13_24, w_stg_0_13_25, w_stg_0_13_26, w_stg_0_13_27, w_stg_0_13_28, w_stg_0_13_29, w_stg_0_13_30, w_stg_0_13_31, w_stg_0_13_32, w_stg_0_13_33, w_stg_0_13_34, w_stg_0_13_35, w_stg_0_13_36, w_stg_0_13_37, w_stg_0_13_38, w_stg_0_13_39, w_stg_0_13_40, w_stg_0_13_41, w_stg_0_13_42, w_stg_0_13_43, w_stg_0_13_44, w_stg_0_14_14, w_stg_0_14_15, w_stg_0_14_16, w_stg_0_14_17, w_stg_0_14_18, w_stg_0_14_19, w_stg_0_14_20, w_stg_0_14_21, w_stg_0_14_22, w_stg_0_14_23, w_stg_0_14_24, w_stg_0_14_25, w_stg_0_14_26, w_stg_0_14_27, w_stg_0_14_28, w_stg_0_14_29, w_stg_0_14_30, w_stg_0_14_31, w_stg_0_14_32, w_stg_0_14_33, w_stg_0_14_34, w_stg_0_14_35, w_stg_0_14_36, w_stg_0_14_37, w_stg_0_14_38, w_stg_0_14_39, w_stg_0_14_40, w_stg_0_14_41, w_stg_0_14_42, w_stg_0_14_43, w_stg_0_14_44, w_stg_0_14_45, w_stg_0_15_15, w_stg_0_15_16, w_stg_0_15_17, w_stg_0_15_18, w_stg_0_15_19, w_stg_0_15_20, w_stg_0_15_21, w_stg_0_15_22, w_stg_0_15_23, w_stg_0_15_24, w_stg_0_15_25, w_stg_0_15_26, w_stg_0_15_27, w_stg_0_15_28, w_stg_0_15_29, w_stg_0_15_30, w_stg_0_15_31, w_stg_0_15_32, w_stg_0_15_33, w_stg_0_15_34, w_stg_0_15_35, w_stg_0_15_36, w_stg_0_15_37, w_stg_0_15_38, w_stg_0_15_39, w_stg_0_15_40, w_stg_0_15_41, w_stg_0_15_42, w_stg_0_15_43, w_stg_0_15_44, w_stg_0_15_45, w_stg_0_15_46, w_stg_0_16_16, w_stg_0_16_17, w_stg_0_16_18, w_stg_0_16_19, w_stg_0_16_20, w_stg_0_16_21, w_stg_0_16_22, w_stg_0_16_23, w_stg_0_16_24, w_stg_0_16_25, w_stg_0_16_26, w_stg_0_16_27, w_stg_0_16_28, w_stg_0_16_29, w_stg_0_16_30, w_stg_0_16_31, w_stg_0_16_32, w_stg_0_16_33, w_stg_0_16_34, w_stg_0_16_35, w_stg_0_16_36, w_stg_0_16_37, w_stg_0_16_38, w_stg_0_16_39, w_stg_0_16_40, w_stg_0_16_41, w_stg_0_16_42, w_stg_0_16_43, w_stg_0_16_44, w_stg_0_16_45, w_stg_0_16_46, w_stg_0_16_47, w_stg_0_17_17, w_stg_0_17_18, w_stg_0_17_19, w_stg_0_17_20, w_stg_0_17_21, w_stg_0_17_22, w_stg_0_17_23, w_stg_0_17_24, w_stg_0_17_25, w_stg_0_17_26, w_stg_0_17_27, w_stg_0_17_28, w_stg_0_17_29, w_stg_0_17_30, w_stg_0_17_31, w_stg_0_17_32, w_stg_0_17_33, w_stg_0_17_34, w_stg_0_17_35, w_stg_0_17_36, w_stg_0_17_37, w_stg_0_17_38, w_stg_0_17_39, w_stg_0_17_40, w_stg_0_17_41, w_stg_0_17_42, w_stg_0_17_43, w_stg_0_17_44, w_stg_0_17_45, w_stg_0_17_46, w_stg_0_17_47, w_stg_0_17_48, w_stg_0_18_18, w_stg_0_18_19, w_stg_0_18_20, w_stg_0_18_21, w_stg_0_18_22, w_stg_0_18_23, w_stg_0_18_24, w_stg_0_18_25, w_stg_0_18_26, w_stg_0_18_27, w_stg_0_18_28, w_stg_0_18_29, w_stg_0_18_30, w_stg_0_18_31, w_stg_0_18_32, w_stg_0_18_33, w_stg_0_18_34, w_stg_0_18_35, w_stg_0_18_36, w_stg_0_18_37, w_stg_0_18_38, w_stg_0_18_39, w_stg_0_18_40, w_stg_0_18_41, w_stg_0_18_42, w_stg_0_18_43, w_stg_0_18_44, w_stg_0_18_45, w_stg_0_18_46, w_stg_0_18_47, w_stg_0_18_48, w_stg_0_18_49, w_stg_0_19_19, w_stg_0_19_20, w_stg_0_19_21, w_stg_0_19_22, w_stg_0_19_23, w_stg_0_19_24, w_stg_0_19_25, w_stg_0_19_26, w_stg_0_19_27, w_stg_0_19_28, w_stg_0_19_29, w_stg_0_19_30, w_stg_0_19_31, w_stg_0_19_32, w_stg_0_19_33, w_stg_0_19_34, w_stg_0_19_35, w_stg_0_19_36, w_stg_0_19_37, w_stg_0_19_38, w_stg_0_19_39, w_stg_0_19_40, w_stg_0_19_41, w_stg_0_19_42, w_stg_0_19_43, w_stg_0_19_44, w_stg_0_19_45, w_stg_0_19_46, w_stg_0_19_47, w_stg_0_19_48, w_stg_0_19_49, w_stg_0_19_50, w_stg_0_20_20, w_stg_0_20_21, w_stg_0_20_22, w_stg_0_20_23, w_stg_0_20_24, w_stg_0_20_25, w_stg_0_20_26, w_stg_0_20_27, w_stg_0_20_28, w_stg_0_20_29, w_stg_0_20_30, w_stg_0_20_31, w_stg_0_20_32, w_stg_0_20_33, w_stg_0_20_34, w_stg_0_20_35, w_stg_0_20_36, w_stg_0_20_37, w_stg_0_20_38, w_stg_0_20_39, w_stg_0_20_40, w_stg_0_20_41, w_stg_0_20_42, w_stg_0_20_43, w_stg_0_20_44, w_stg_0_20_45, w_stg_0_20_46, w_stg_0_20_47, w_stg_0_20_48, w_stg_0_20_49, w_stg_0_20_50, w_stg_0_20_51, w_stg_0_21_21, w_stg_0_21_22, w_stg_0_21_23, w_stg_0_21_24, w_stg_0_21_25, w_stg_0_21_26, w_stg_0_21_27, w_stg_0_21_28, w_stg_0_21_29, w_stg_0_21_30, w_stg_0_21_31, w_stg_0_21_32, w_stg_0_21_33, w_stg_0_21_34, w_stg_0_21_35, w_stg_0_21_36, w_stg_0_21_37, w_stg_0_21_38, w_stg_0_21_39, w_stg_0_21_40, w_stg_0_21_41, w_stg_0_21_42, w_stg_0_21_43, w_stg_0_21_44, w_stg_0_21_45, w_stg_0_21_46, w_stg_0_21_47, w_stg_0_21_48, w_stg_0_21_49, w_stg_0_21_50, w_stg_0_21_51, w_stg_0_21_52, w_stg_0_22_22, w_stg_0_22_23, w_stg_0_22_24, w_stg_0_22_25, w_stg_0_22_26, w_stg_0_22_27, w_stg_0_22_28, w_stg_0_22_29, w_stg_0_22_30, w_stg_0_22_31, w_stg_0_22_32, w_stg_0_22_33, w_stg_0_22_34, w_stg_0_22_35, w_stg_0_22_36, w_stg_0_22_37, w_stg_0_22_38, w_stg_0_22_39, w_stg_0_22_40, w_stg_0_22_41, w_stg_0_22_42, w_stg_0_22_43, w_stg_0_22_44, w_stg_0_22_45, w_stg_0_22_46, w_stg_0_22_47, w_stg_0_22_48, w_stg_0_22_49, w_stg_0_22_50, w_stg_0_22_51, w_stg_0_22_52, w_stg_0_22_53, w_stg_0_23_23, w_stg_0_23_24, w_stg_0_23_25, w_stg_0_23_26, w_stg_0_23_27, w_stg_0_23_28, w_stg_0_23_29, w_stg_0_23_30, w_stg_0_23_31, w_stg_0_23_32, w_stg_0_23_33, w_stg_0_23_34, w_stg_0_23_35, w_stg_0_23_36, w_stg_0_23_37, w_stg_0_23_38, w_stg_0_23_39, w_stg_0_23_40, w_stg_0_23_41, w_stg_0_23_42, w_stg_0_23_43, w_stg_0_23_44, w_stg_0_23_45, w_stg_0_23_46, w_stg_0_23_47, w_stg_0_23_48, w_stg_0_23_49, w_stg_0_23_50, w_stg_0_23_51, w_stg_0_23_52, w_stg_0_23_53, w_stg_0_23_54, w_stg_0_24_24, w_stg_0_24_25, w_stg_0_24_26, w_stg_0_24_27, w_stg_0_24_28, w_stg_0_24_29, w_stg_0_24_30, w_stg_0_24_31, w_stg_0_24_32, w_stg_0_24_33, w_stg_0_24_34, w_stg_0_24_35, w_stg_0_24_36, w_stg_0_24_37, w_stg_0_24_38, w_stg_0_24_39, w_stg_0_24_40, w_stg_0_24_41, w_stg_0_24_42, w_stg_0_24_43, w_stg_0_24_44, w_stg_0_24_45, w_stg_0_24_46, w_stg_0_24_47, w_stg_0_24_48, w_stg_0_24_49, w_stg_0_24_50, w_stg_0_24_51, w_stg_0_24_52, w_stg_0_24_53, w_stg_0_24_54, w_stg_0_24_55, w_stg_0_25_25, w_stg_0_25_26, w_stg_0_25_27, w_stg_0_25_28, w_stg_0_25_29, w_stg_0_25_30, w_stg_0_25_31, w_stg_0_25_32, w_stg_0_25_33, w_stg_0_25_34, w_stg_0_25_35, w_stg_0_25_36, w_stg_0_25_37, w_stg_0_25_38, w_stg_0_25_39, w_stg_0_25_40, w_stg_0_25_41, w_stg_0_25_42, w_stg_0_25_43, w_stg_0_25_44, w_stg_0_25_45, w_stg_0_25_46, w_stg_0_25_47, w_stg_0_25_48, w_stg_0_25_49, w_stg_0_25_50, w_stg_0_25_51, w_stg_0_25_52, w_stg_0_25_53, w_stg_0_25_54, w_stg_0_25_55, w_stg_0_25_56, w_stg_0_26_26, w_stg_0_26_27, w_stg_0_26_28, w_stg_0_26_29, w_stg_0_26_30, w_stg_0_26_31, w_stg_0_26_32, w_stg_0_26_33, w_stg_0_26_34, w_stg_0_26_35, w_stg_0_26_36, w_stg_0_26_37, w_stg_0_26_38, w_stg_0_26_39, w_stg_0_26_40, w_stg_0_26_41, w_stg_0_26_42, w_stg_0_26_43, w_stg_0_26_44, w_stg_0_26_45, w_stg_0_26_46, w_stg_0_26_47, w_stg_0_26_48, w_stg_0_26_49, w_stg_0_26_50, w_stg_0_26_51, w_stg_0_26_52, w_stg_0_26_53, w_stg_0_26_54, w_stg_0_26_55, w_stg_0_26_56, w_stg_0_26_57, w_stg_0_27_27, w_stg_0_27_28, w_stg_0_27_29, w_stg_0_27_30, w_stg_0_27_31, w_stg_0_27_32, w_stg_0_27_33, w_stg_0_27_34, w_stg_0_27_35, w_stg_0_27_36, w_stg_0_27_37, w_stg_0_27_38, w_stg_0_27_39, w_stg_0_27_40, w_stg_0_27_41, w_stg_0_27_42, w_stg_0_27_43, w_stg_0_27_44, w_stg_0_27_45, w_stg_0_27_46, w_stg_0_27_47, w_stg_0_27_48, w_stg_0_27_49, w_stg_0_27_50, w_stg_0_27_51, w_stg_0_27_52, w_stg_0_27_53, w_stg_0_27_54, w_stg_0_27_55, w_stg_0_27_56, w_stg_0_27_57, w_stg_0_27_58, w_stg_0_28_28, w_stg_0_28_29, w_stg_0_28_30, w_stg_0_28_31, w_stg_0_28_32, w_stg_0_28_33, w_stg_0_28_34, w_stg_0_28_35, w_stg_0_28_36, w_stg_0_28_37, w_stg_0_28_38, w_stg_0_28_39, w_stg_0_28_40, w_stg_0_28_41, w_stg_0_28_42, w_stg_0_28_43, w_stg_0_28_44, w_stg_0_28_45, w_stg_0_28_46, w_stg_0_28_47, w_stg_0_28_48, w_stg_0_28_49, w_stg_0_28_50, w_stg_0_28_51, w_stg_0_28_52, w_stg_0_28_53, w_stg_0_28_54, w_stg_0_28_55, w_stg_0_28_56, w_stg_0_28_57, w_stg_0_28_58, w_stg_0_28_59, w_stg_0_29_29, w_stg_0_29_30, w_stg_0_29_31, w_stg_0_29_32, w_stg_0_29_33, w_stg_0_29_34, w_stg_0_29_35, w_stg_0_29_36, w_stg_0_29_37, w_stg_0_29_38, w_stg_0_29_39, w_stg_0_29_40, w_stg_0_29_41, w_stg_0_29_42, w_stg_0_29_43, w_stg_0_29_44, w_stg_0_29_45, w_stg_0_29_46, w_stg_0_29_47, w_stg_0_29_48, w_stg_0_29_49, w_stg_0_29_50, w_stg_0_29_51, w_stg_0_29_52, w_stg_0_29_53, w_stg_0_29_54, w_stg_0_29_55, w_stg_0_29_56, w_stg_0_29_57, w_stg_0_29_58, w_stg_0_29_59, w_stg_0_29_60, w_stg_0_30_30, w_stg_0_30_31, w_stg_0_30_32, w_stg_0_30_33, w_stg_0_30_34, w_stg_0_30_35, w_stg_0_30_36, w_stg_0_30_37, w_stg_0_30_38, w_stg_0_30_39, w_stg_0_30_40, w_stg_0_30_41, w_stg_0_30_42, w_stg_0_30_43, w_stg_0_30_44, w_stg_0_30_45, w_stg_0_30_46, w_stg_0_30_47, w_stg_0_30_48, w_stg_0_30_49, w_stg_0_30_50, w_stg_0_30_51, w_stg_0_30_52, w_stg_0_30_53, w_stg_0_30_54, w_stg_0_30_55, w_stg_0_30_56, w_stg_0_30_57, w_stg_0_30_58, w_stg_0_30_59, w_stg_0_30_60, w_stg_0_30_61, w_stg_0_31_31, w_stg_0_31_32, w_stg_0_31_33, w_stg_0_31_34, w_stg_0_31_35, w_stg_0_31_36, w_stg_0_31_37, w_stg_0_31_38, w_stg_0_31_39, w_stg_0_31_40, w_stg_0_31_41, w_stg_0_31_42, w_stg_0_31_43, w_stg_0_31_44, w_stg_0_31_45, w_stg_0_31_46, w_stg_0_31_47, w_stg_0_31_48, w_stg_0_31_49, w_stg_0_31_50, w_stg_0_31_51, w_stg_0_31_52, w_stg_0_31_53, w_stg_0_31_54, w_stg_0_31_55, w_stg_0_31_56, w_stg_0_31_57, w_stg_0_31_58, w_stg_0_31_59, w_stg_0_31_60, w_stg_0_31_61, w_stg_0_31_62;
	wire w_stg_1_0_0, w_stg_1_0_1, w_stg_1_0_2, w_stg_1_1_2, w_stg_1_0_3, w_stg_1_1_3, w_stg_1_0_4, w_stg_1_2_3, w_stg_1_1_4, w_stg_1_0_5, w_stg_1_2_4, w_stg_1_1_5, w_stg_1_2_5, w_stg_1_0_6, w_stg_1_3_5, w_stg_1_1_6, w_stg_1_2_6, w_stg_1_0_7, w_stg_1_3_6, w_stg_1_1_7, w_stg_1_4_6, w_stg_1_2_7, w_stg_1_0_8, w_stg_1_3_7, w_stg_1_1_8, w_stg_1_4_7, w_stg_1_2_8, w_stg_1_3_8, w_stg_1_0_9, w_stg_1_4_8, w_stg_1_1_9, w_stg_1_5_8, w_stg_1_2_9, w_stg_1_3_9, w_stg_1_0_10, w_stg_1_4_9, w_stg_1_1_10, w_stg_1_5_9, w_stg_1_2_10, w_stg_1_6_9, w_stg_1_3_10, w_stg_1_0_11, w_stg_1_4_10, w_stg_1_1_11, w_stg_1_5_10, w_stg_1_2_11, w_stg_1_6_10, w_stg_1_3_11, w_stg_1_4_11, w_stg_1_0_12, w_stg_1_5_11, w_stg_1_1_12, w_stg_1_6_11, w_stg_1_2_12, w_stg_1_7_11, w_stg_1_3_12, w_stg_1_4_12, w_stg_1_0_13, w_stg_1_5_12, w_stg_1_1_13, w_stg_1_6_12, w_stg_1_2_13, w_stg_1_7_12, w_stg_1_3_13, w_stg_1_8_12, w_stg_1_4_13, w_stg_1_0_14, w_stg_1_5_13, w_stg_1_1_14, w_stg_1_6_13, w_stg_1_2_14, w_stg_1_7_13, w_stg_1_3_14, w_stg_1_8_13, w_stg_1_4_14, w_stg_1_5_14, w_stg_1_0_15, w_stg_1_6_14, w_stg_1_1_15, w_stg_1_7_14, w_stg_1_2_15, w_stg_1_8_14, w_stg_1_3_15, w_stg_1_9_14, w_stg_1_4_15, w_stg_1_5_15, w_stg_1_0_16, w_stg_1_6_15, w_stg_1_1_16, w_stg_1_7_15, w_stg_1_2_16, w_stg_1_8_15, w_stg_1_3_16, w_stg_1_9_15, w_stg_1_4_16, w_stg_1_10_15, w_stg_1_5_16, w_stg_1_0_17, w_stg_1_6_16, w_stg_1_1_17, w_stg_1_7_16, w_stg_1_2_17, w_stg_1_8_16, w_stg_1_3_17, w_stg_1_9_16, w_stg_1_4_17, w_stg_1_10_16, w_stg_1_5_17, w_stg_1_6_17, w_stg_1_0_18, w_stg_1_7_17, w_stg_1_1_18, w_stg_1_8_17, w_stg_1_2_18, w_stg_1_9_17, w_stg_1_3_18, w_stg_1_10_17, w_stg_1_4_18, w_stg_1_11_17, w_stg_1_5_18, w_stg_1_6_18, w_stg_1_0_19, w_stg_1_7_18, w_stg_1_1_19, w_stg_1_8_18, w_stg_1_2_19, w_stg_1_9_18, w_stg_1_3_19, w_stg_1_10_18, w_stg_1_4_19, w_stg_1_11_18, w_stg_1_5_19, w_stg_1_12_18, w_stg_1_6_19, w_stg_1_0_20, w_stg_1_7_19, w_stg_1_1_20, w_stg_1_8_19, w_stg_1_2_20, w_stg_1_9_19, w_stg_1_3_20, w_stg_1_10_19, w_stg_1_4_20, w_stg_1_11_19, w_stg_1_5_20, w_stg_1_12_19, w_stg_1_6_20, w_stg_1_7_20, w_stg_1_0_21, w_stg_1_8_20, w_stg_1_1_21, w_stg_1_9_20, w_stg_1_2_21, w_stg_1_10_20, w_stg_1_3_21, w_stg_1_11_20, w_stg_1_4_21, w_stg_1_12_20, w_stg_1_5_21, w_stg_1_13_20, w_stg_1_6_21, w_stg_1_7_21, w_stg_1_0_22, w_stg_1_8_21, w_stg_1_1_22, w_stg_1_9_21, w_stg_1_2_22, w_stg_1_10_21, w_stg_1_3_22, w_stg_1_11_21, w_stg_1_4_22, w_stg_1_12_21, w_stg_1_5_22, w_stg_1_13_21, w_stg_1_6_22, w_stg_1_14_21, w_stg_1_7_22, w_stg_1_0_23, w_stg_1_8_22, w_stg_1_1_23, w_stg_1_9_22, w_stg_1_2_23, w_stg_1_10_22, w_stg_1_3_23, w_stg_1_11_22, w_stg_1_4_23, w_stg_1_12_22, w_stg_1_5_23, w_stg_1_13_22, w_stg_1_6_23, w_stg_1_14_22, w_stg_1_7_23, w_stg_1_8_23, w_stg_1_0_24, w_stg_1_9_23, w_stg_1_1_24, w_stg_1_10_23, w_stg_1_2_24, w_stg_1_11_23, w_stg_1_3_24, w_stg_1_12_23, w_stg_1_4_24, w_stg_1_13_23, w_stg_1_5_24, w_stg_1_14_23, w_stg_1_6_24, w_stg_1_15_23, w_stg_1_7_24, w_stg_1_8_24, w_stg_1_0_25, w_stg_1_9_24, w_stg_1_1_25, w_stg_1_10_24, w_stg_1_2_25, w_stg_1_11_24, w_stg_1_3_25, w_stg_1_12_24, w_stg_1_4_25, w_stg_1_13_24, w_stg_1_5_25, w_stg_1_14_24, w_stg_1_6_25, w_stg_1_15_24, w_stg_1_7_25, w_stg_1_16_24, w_stg_1_8_25, w_stg_1_0_26, w_stg_1_9_25, w_stg_1_1_26, w_stg_1_10_25, w_stg_1_2_26, w_stg_1_11_25, w_stg_1_3_26, w_stg_1_12_25, w_stg_1_4_26, w_stg_1_13_25, w_stg_1_5_26, w_stg_1_14_25, w_stg_1_6_26, w_stg_1_15_25, w_stg_1_7_26, w_stg_1_16_25, w_stg_1_8_26, w_stg_1_9_26, w_stg_1_0_27, w_stg_1_10_26, w_stg_1_1_27, w_stg_1_11_26, w_stg_1_2_27, w_stg_1_12_26, w_stg_1_3_27, w_stg_1_13_26, w_stg_1_4_27, w_stg_1_14_26, w_stg_1_5_27, w_stg_1_15_26, w_stg_1_6_27, w_stg_1_16_26, w_stg_1_7_27, w_stg_1_17_26, w_stg_1_8_27, w_stg_1_9_27, w_stg_1_0_28, w_stg_1_10_27, w_stg_1_1_28, w_stg_1_11_27, w_stg_1_2_28, w_stg_1_12_27, w_stg_1_3_28, w_stg_1_13_27, w_stg_1_4_28, w_stg_1_14_27, w_stg_1_5_28, w_stg_1_15_27, w_stg_1_6_28, w_stg_1_16_27, w_stg_1_7_28, w_stg_1_17_27, w_stg_1_8_28, w_stg_1_18_27, w_stg_1_9_28, w_stg_1_0_29, w_stg_1_10_28, w_stg_1_1_29, w_stg_1_11_28, w_stg_1_2_29, w_stg_1_12_28, w_stg_1_3_29, w_stg_1_13_28, w_stg_1_4_29, w_stg_1_14_28, w_stg_1_5_29, w_stg_1_15_28, w_stg_1_6_29, w_stg_1_16_28, w_stg_1_7_29, w_stg_1_17_28, w_stg_1_8_29, w_stg_1_18_28, w_stg_1_9_29, w_stg_1_10_29, w_stg_1_0_30, w_stg_1_11_29, w_stg_1_1_30, w_stg_1_12_29, w_stg_1_2_30, w_stg_1_13_29, w_stg_1_3_30, w_stg_1_14_29, w_stg_1_4_30, w_stg_1_15_29, w_stg_1_5_30, w_stg_1_16_29, w_stg_1_6_30, w_stg_1_17_29, w_stg_1_7_30, w_stg_1_18_29, w_stg_1_8_30, w_stg_1_19_29, w_stg_1_9_30, w_stg_1_10_30, w_stg_1_0_31, w_stg_1_11_30, w_stg_1_1_31, w_stg_1_12_30, w_stg_1_2_31, w_stg_1_13_30, w_stg_1_3_31, w_stg_1_14_30, w_stg_1_4_31, w_stg_1_15_30, w_stg_1_5_31, w_stg_1_16_30, w_stg_1_6_31, w_stg_1_17_30, w_stg_1_7_31, w_stg_1_18_30, w_stg_1_8_31, w_stg_1_19_30, w_stg_1_9_31, w_stg_1_20_30, w_stg_1_10_31, w_stg_1_0_32, w_stg_1_11_31, w_stg_1_1_32, w_stg_1_12_31, w_stg_1_2_32, w_stg_1_13_31, w_stg_1_3_32, w_stg_1_14_31, w_stg_1_4_32, w_stg_1_15_31, w_stg_1_5_32, w_stg_1_16_31, w_stg_1_6_32, w_stg_1_17_31, w_stg_1_7_32, w_stg_1_18_31, w_stg_1_8_32, w_stg_1_19_31, w_stg_1_9_32, w_stg_1_20_31, w_stg_1_10_32, w_stg_1_11_32, w_stg_1_0_33, w_stg_1_12_32, w_stg_1_1_33, w_stg_1_13_32, w_stg_1_2_33, w_stg_1_14_32, w_stg_1_3_33, w_stg_1_15_32, w_stg_1_4_33, w_stg_1_16_32, w_stg_1_5_33, w_stg_1_17_32, w_stg_1_6_33, w_stg_1_18_32, w_stg_1_7_33, w_stg_1_19_32, w_stg_1_8_33, w_stg_1_20_32, w_stg_1_9_33, w_stg_1_21_32, w_stg_1_10_33, w_stg_1_11_33, w_stg_1_12_33, w_stg_1_0_34, w_stg_1_13_33, w_stg_1_1_34, w_stg_1_14_33, w_stg_1_2_34, w_stg_1_15_33, w_stg_1_3_34, w_stg_1_16_33, w_stg_1_4_34, w_stg_1_17_33, w_stg_1_5_34, w_stg_1_18_33, w_stg_1_6_34, w_stg_1_19_33, w_stg_1_7_34, w_stg_1_20_33, w_stg_1_8_34, w_stg_1_21_33, w_stg_1_9_34, w_stg_1_10_34, w_stg_1_0_35, w_stg_1_11_34, w_stg_1_1_35, w_stg_1_12_34, w_stg_1_2_35, w_stg_1_13_34, w_stg_1_3_35, w_stg_1_14_34, w_stg_1_4_35, w_stg_1_15_34, w_stg_1_5_35, w_stg_1_16_34, w_stg_1_6_35, w_stg_1_17_34, w_stg_1_7_35, w_stg_1_18_34, w_stg_1_8_35, w_stg_1_19_34, w_stg_1_9_35, w_stg_1_10_35, w_stg_1_0_36, w_stg_1_11_35, w_stg_1_1_36, w_stg_1_12_35, w_stg_1_2_36, w_stg_1_13_35, w_stg_1_3_36, w_stg_1_14_35, w_stg_1_4_36, w_stg_1_15_35, w_stg_1_5_36, w_stg_1_16_35, w_stg_1_6_36, w_stg_1_17_35, w_stg_1_7_36, w_stg_1_18_35, w_stg_1_8_36, w_stg_1_19_35, w_stg_1_9_36, w_stg_1_10_36, w_stg_1_11_36, w_stg_1_0_37, w_stg_1_12_36, w_stg_1_1_37, w_stg_1_13_36, w_stg_1_2_37, w_stg_1_14_36, w_stg_1_3_37, w_stg_1_15_36, w_stg_1_4_37, w_stg_1_16_36, w_stg_1_5_37, w_stg_1_17_36, w_stg_1_6_37, w_stg_1_18_36, w_stg_1_7_37, w_stg_1_19_36, w_stg_1_8_37, w_stg_1_9_37, w_stg_1_0_38, w_stg_1_10_37, w_stg_1_1_38, w_stg_1_11_37, w_stg_1_2_38, w_stg_1_12_37, w_stg_1_3_38, w_stg_1_13_37, w_stg_1_4_38, w_stg_1_14_37, w_stg_1_5_38, w_stg_1_15_37, w_stg_1_6_38, w_stg_1_16_37, w_stg_1_7_38, w_stg_1_17_37, w_stg_1_8_38, w_stg_1_9_38, w_stg_1_0_39, w_stg_1_10_38, w_stg_1_1_39, w_stg_1_11_38, w_stg_1_2_39, w_stg_1_12_38, w_stg_1_3_39, w_stg_1_13_38, w_stg_1_4_39, w_stg_1_14_38, w_stg_1_5_39, w_stg_1_15_38, w_stg_1_6_39, w_stg_1_16_38, w_stg_1_7_39, w_stg_1_17_38, w_stg_1_8_39, w_stg_1_9_39, w_stg_1_10_39, w_stg_1_0_40, w_stg_1_11_39, w_stg_1_1_40, w_stg_1_12_39, w_stg_1_2_40, w_stg_1_13_39, w_stg_1_3_40, w_stg_1_14_39, w_stg_1_4_40, w_stg_1_15_39, w_stg_1_5_40, w_stg_1_16_39, w_stg_1_6_40, w_stg_1_17_39, w_stg_1_7_40, w_stg_1_8_40, w_stg_1_0_41, w_stg_1_9_40, w_stg_1_1_41, w_stg_1_10_40, w_stg_1_2_41, w_stg_1_11_40, w_stg_1_3_41, w_stg_1_12_40, w_stg_1_4_41, w_stg_1_13_40, w_stg_1_5_41, w_stg_1_14_40, w_stg_1_6_41, w_stg_1_15_40, w_stg_1_7_41, w_stg_1_8_41, w_stg_1_0_42, w_stg_1_9_41, w_stg_1_1_42, w_stg_1_10_41, w_stg_1_2_42, w_stg_1_11_41, w_stg_1_3_42, w_stg_1_12_41, w_stg_1_4_42, w_stg_1_13_41, w_stg_1_5_42, w_stg_1_14_41, w_stg_1_6_42, w_stg_1_15_41, w_stg_1_7_42, w_stg_1_8_42, w_stg_1_9_42, w_stg_1_0_43, w_stg_1_10_42, w_stg_1_1_43, w_stg_1_11_42, w_stg_1_2_43, w_stg_1_12_42, w_stg_1_3_43, w_stg_1_13_42, w_stg_1_4_43, w_stg_1_14_42, w_stg_1_5_43, w_stg_1_15_42, w_stg_1_6_43, w_stg_1_7_43, w_stg_1_0_44, w_stg_1_8_43, w_stg_1_1_44, w_stg_1_9_43, w_stg_1_2_44, w_stg_1_10_43, w_stg_1_3_44, w_stg_1_11_43, w_stg_1_4_44, w_stg_1_12_43, w_stg_1_5_44, w_stg_1_13_43, w_stg_1_6_44, w_stg_1_7_44, w_stg_1_0_45, w_stg_1_8_44, w_stg_1_1_45, w_stg_1_9_44, w_stg_1_2_45, w_stg_1_10_44, w_stg_1_3_45, w_stg_1_11_44, w_stg_1_4_45, w_stg_1_12_44, w_stg_1_5_45, w_stg_1_13_44, w_stg_1_6_45, w_stg_1_7_45, w_stg_1_8_45, w_stg_1_0_46, w_stg_1_9_45, w_stg_1_1_46, w_stg_1_10_45, w_stg_1_2_46, w_stg_1_11_45, w_stg_1_3_46, w_stg_1_12_45, w_stg_1_4_46, w_stg_1_13_45, w_stg_1_5_46, w_stg_1_6_46, w_stg_1_0_47, w_stg_1_7_46, w_stg_1_1_47, w_stg_1_8_46, w_stg_1_2_47, w_stg_1_9_46, w_stg_1_3_47, w_stg_1_10_46, w_stg_1_4_47, w_stg_1_11_46, w_stg_1_5_47, w_stg_1_6_47, w_stg_1_0_48, w_stg_1_7_47, w_stg_1_1_48, w_stg_1_8_47, w_stg_1_2_48, w_stg_1_9_47, w_stg_1_3_48, w_stg_1_10_47, w_stg_1_4_48, w_stg_1_11_47, w_stg_1_5_48, w_stg_1_6_48, w_stg_1_7_48, w_stg_1_0_49, w_stg_1_8_48, w_stg_1_1_49, w_stg_1_9_48, w_stg_1_2_49, w_stg_1_10_48, w_stg_1_3_49, w_stg_1_11_48, w_stg_1_4_49, w_stg_1_5_49, w_stg_1_0_50, w_stg_1_6_49, w_stg_1_1_50, w_stg_1_7_49, w_stg_1_2_50, w_stg_1_8_49, w_stg_1_3_50, w_stg_1_9_49, w_stg_1_4_50, w_stg_1_5_50, w_stg_1_0_51, w_stg_1_6_50, w_stg_1_1_51, w_stg_1_7_50, w_stg_1_2_51, w_stg_1_8_50, w_stg_1_3_51, w_stg_1_9_50, w_stg_1_4_51, w_stg_1_5_51, w_stg_1_6_51, w_stg_1_0_52, w_stg_1_7_51, w_stg_1_1_52, w_stg_1_8_51, w_stg_1_2_52, w_stg_1_9_51, w_stg_1_3_52, w_stg_1_4_52, w_stg_1_0_53, w_stg_1_5_52, w_stg_1_1_53, w_stg_1_6_52, w_stg_1_2_53, w_stg_1_7_52, w_stg_1_3_53, w_stg_1_4_53, w_stg_1_0_54, w_stg_1_5_53, w_stg_1_1_54, w_stg_1_6_53, w_stg_1_2_54, w_stg_1_7_53, w_stg_1_3_54, w_stg_1_4_54, w_stg_1_5_54, w_stg_1_0_55, w_stg_1_6_54, w_stg_1_1_55, w_stg_1_7_54, w_stg_1_2_55, w_stg_1_3_55, w_stg_1_0_56, w_stg_1_4_55, w_stg_1_1_56, w_stg_1_5_55, w_stg_1_2_56, w_stg_1_3_56, w_stg_1_0_57, w_stg_1_4_56, w_stg_1_1_57, w_stg_1_5_56, w_stg_1_2_57, w_stg_1_3_57, w_stg_1_4_57, w_stg_1_0_58, w_stg_1_5_57, w_stg_1_1_58, w_stg_1_2_58, w_stg_1_0_59, w_stg_1_3_58, w_stg_1_1_59, w_stg_1_2_59, w_stg_1_0_60, w_stg_1_3_59, w_stg_1_1_60, w_stg_1_2_60, w_stg_1_3_60, w_stg_1_0_61, w_stg_1_1_61, w_stg_1_0_62, w_stg_1_1_62;
	wire w_stg_2_0_0, w_stg_2_0_1, w_stg_2_0_2, w_stg_2_0_3, w_stg_2_1_3, w_stg_2_0_4, w_stg_2_1_4, w_stg_2_0_5, w_stg_2_1_5, w_stg_2_0_6, w_stg_2_2_5, w_stg_2_1_6, w_stg_2_0_7, w_stg_2_2_6, w_stg_2_1_7, w_stg_2_2_7, w_stg_2_0_8, w_stg_2_3_7, w_stg_2_1_8, w_stg_2_2_8, w_stg_2_0_9, w_stg_2_3_8, w_stg_2_1_9, w_stg_2_2_9, w_stg_2_0_10, w_stg_2_3_9, w_stg_2_1_10, w_stg_2_4_9, w_stg_2_2_10, w_stg_2_0_11, w_stg_2_3_10, w_stg_2_1_11, w_stg_2_4_10, w_stg_2_2_11, w_stg_2_0_12, w_stg_2_3_11, w_stg_2_1_12, w_stg_2_4_11, w_stg_2_2_12, w_stg_2_3_12, w_stg_2_0_13, w_stg_2_4_12, w_stg_2_1_13, w_stg_2_5_12, w_stg_2_2_13, w_stg_2_3_13, w_stg_2_0_14, w_stg_2_4_13, w_stg_2_1_14, w_stg_2_5_13, w_stg_2_2_14, w_stg_2_3_14, w_stg_2_0_15, w_stg_2_4_14, w_stg_2_1_15, w_stg_2_5_14, w_stg_2_2_15, w_stg_2_6_14, w_stg_2_3_15, w_stg_2_0_16, w_stg_2_4_15, w_stg_2_1_16, w_stg_2_5_15, w_stg_2_2_16, w_stg_2_6_15, w_stg_2_3_16, w_stg_2_4_16, w_stg_2_0_17, w_stg_2_5_16, w_stg_2_1_17, w_stg_2_6_16, w_stg_2_2_17, w_stg_2_7_16, w_stg_2_3_17, w_stg_2_4_17, w_stg_2_0_18, w_stg_2_5_17, w_stg_2_1_18, w_stg_2_6_17, w_stg_2_2_18, w_stg_2_7_17, w_stg_2_3_18, w_stg_2_4_18, w_stg_2_0_19, w_stg_2_5_18, w_stg_2_1_19, w_stg_2_6_18, w_stg_2_2_19, w_stg_2_7_18, w_stg_2_3_19, w_stg_2_8_18, w_stg_2_4_19, w_stg_2_0_20, w_stg_2_5_19, w_stg_2_1_20, w_stg_2_6_19, w_stg_2_2_20, w_stg_2_7_19, w_stg_2_3_20, w_stg_2_8_19, w_stg_2_4_20, w_stg_2_0_21, w_stg_2_5_20, w_stg_2_1_21, w_stg_2_6_20, w_stg_2_2_21, w_stg_2_7_20, w_stg_2_3_21, w_stg_2_8_20, w_stg_2_4_21, w_stg_2_5_21, w_stg_2_0_22, w_stg_2_6_21, w_stg_2_1_22, w_stg_2_7_21, w_stg_2_2_22, w_stg_2_8_21, w_stg_2_3_22, w_stg_2_9_21, w_stg_2_4_22, w_stg_2_5_22, w_stg_2_0_23, w_stg_2_6_22, w_stg_2_1_23, w_stg_2_7_22, w_stg_2_2_23, w_stg_2_8_22, w_stg_2_3_23, w_stg_2_9_22, w_stg_2_4_23, w_stg_2_5_23, w_stg_2_0_24, w_stg_2_6_23, w_stg_2_1_24, w_stg_2_7_23, w_stg_2_2_24, w_stg_2_8_23, w_stg_2_3_24, w_stg_2_9_23, w_stg_2_4_24, w_stg_2_10_23, w_stg_2_5_24, w_stg_2_0_25, w_stg_2_6_24, w_stg_2_1_25, w_stg_2_7_24, w_stg_2_2_25, w_stg_2_8_24, w_stg_2_3_25, w_stg_2_9_24, w_stg_2_4_25, w_stg_2_10_24, w_stg_2_5_25, w_stg_2_6_25, w_stg_2_0_26, w_stg_2_7_25, w_stg_2_1_26, w_stg_2_8_25, w_stg_2_2_26, w_stg_2_9_25, w_stg_2_3_26, w_stg_2_10_25, w_stg_2_4_26, w_stg_2_11_25, w_stg_2_5_26, w_stg_2_6_26, w_stg_2_0_27, w_stg_2_7_26, w_stg_2_1_27, w_stg_2_8_26, w_stg_2_2_27, w_stg_2_9_26, w_stg_2_3_27, w_stg_2_10_26, w_stg_2_4_27, w_stg_2_11_26, w_stg_2_5_27, w_stg_2_6_27, w_stg_2_0_28, w_stg_2_7_27, w_stg_2_1_28, w_stg_2_8_27, w_stg_2_2_28, w_stg_2_9_27, w_stg_2_3_28, w_stg_2_10_27, w_stg_2_4_28, w_stg_2_11_27, w_stg_2_5_28, w_stg_2_12_27, w_stg_2_6_28, w_stg_2_0_29, w_stg_2_7_28, w_stg_2_1_29, w_stg_2_8_28, w_stg_2_2_29, w_stg_2_9_28, w_stg_2_3_29, w_stg_2_10_28, w_stg_2_4_29, w_stg_2_11_28, w_stg_2_5_29, w_stg_2_12_28, w_stg_2_6_29, w_stg_2_0_30, w_stg_2_7_29, w_stg_2_1_30, w_stg_2_8_29, w_stg_2_2_30, w_stg_2_9_29, w_stg_2_3_30, w_stg_2_10_29, w_stg_2_4_30, w_stg_2_11_29, w_stg_2_5_30, w_stg_2_12_29, w_stg_2_6_30, w_stg_2_7_30, w_stg_2_0_31, w_stg_2_8_30, w_stg_2_1_31, w_stg_2_9_30, w_stg_2_2_31, w_stg_2_10_30, w_stg_2_3_31, w_stg_2_11_30, w_stg_2_4_31, w_stg_2_12_30, w_stg_2_5_31, w_stg_2_13_30, w_stg_2_6_31, w_stg_2_7_31, w_stg_2_0_32, w_stg_2_8_31, w_stg_2_1_32, w_stg_2_9_31, w_stg_2_2_32, w_stg_2_10_31, w_stg_2_3_32, w_stg_2_11_31, w_stg_2_4_32, w_stg_2_12_31, w_stg_2_5_32, w_stg_2_13_31, w_stg_2_6_32, w_stg_2_7_32, w_stg_2_0_33, w_stg_2_8_32, w_stg_2_1_33, w_stg_2_9_32, w_stg_2_2_33, w_stg_2_10_32, w_stg_2_3_33, w_stg_2_11_32, w_stg_2_4_33, w_stg_2_12_32, w_stg_2_5_33, w_stg_2_13_32, w_stg_2_6_33, w_stg_2_14_32, w_stg_2_7_33, w_stg_2_0_34, w_stg_2_8_33, w_stg_2_1_34, w_stg_2_9_33, w_stg_2_2_34, w_stg_2_10_33, w_stg_2_3_34, w_stg_2_11_33, w_stg_2_4_34, w_stg_2_12_33, w_stg_2_5_34, w_stg_2_13_33, w_stg_2_6_34, w_stg_2_14_33, w_stg_2_7_34, w_stg_2_0_35, w_stg_2_8_34, w_stg_2_1_35, w_stg_2_9_34, w_stg_2_2_35, w_stg_2_10_34, w_stg_2_3_35, w_stg_2_11_34, w_stg_2_4_35, w_stg_2_12_34, w_stg_2_5_35, w_stg_2_13_34, w_stg_2_6_35, w_stg_2_7_35, w_stg_2_0_36, w_stg_2_8_35, w_stg_2_1_36, w_stg_2_9_35, w_stg_2_2_36, w_stg_2_10_35, w_stg_2_3_36, w_stg_2_11_35, w_stg_2_4_36, w_stg_2_12_35, w_stg_2_5_36, w_stg_2_13_35, w_stg_2_6_36, w_stg_2_7_36, w_stg_2_0_37, w_stg_2_8_36, w_stg_2_1_37, w_stg_2_9_36, w_stg_2_2_37, w_stg_2_10_36, w_stg_2_3_37, w_stg_2_11_36, w_stg_2_4_37, w_stg_2_12_36, w_stg_2_5_37, w_stg_2_13_36, w_stg_2_6_37, w_stg_2_7_37, w_stg_2_0_38, w_stg_2_8_37, w_stg_2_1_38, w_stg_2_9_37, w_stg_2_2_38, w_stg_2_10_37, w_stg_2_3_38, w_stg_2_11_37, w_stg_2_4_38, w_stg_2_12_37, w_stg_2_5_38, w_stg_2_6_38, w_stg_2_0_39, w_stg_2_7_38, w_stg_2_1_39, w_stg_2_8_38, w_stg_2_2_39, w_stg_2_9_38, w_stg_2_3_39, w_stg_2_10_38, w_stg_2_4_39, w_stg_2_11_38, w_stg_2_5_39, w_stg_2_6_39, w_stg_2_0_40, w_stg_2_7_39, w_stg_2_1_40, w_stg_2_8_39, w_stg_2_2_40, w_stg_2_9_39, w_stg_2_3_40, w_stg_2_10_39, w_stg_2_4_40, w_stg_2_11_39, w_stg_2_5_40, w_stg_2_6_40, w_stg_2_0_41, w_stg_2_7_40, w_stg_2_1_41, w_stg_2_8_40, w_stg_2_2_41, w_stg_2_9_40, w_stg_2_3_41, w_stg_2_10_40, w_stg_2_4_41, w_stg_2_11_40, w_stg_2_5_41, w_stg_2_0_42, w_stg_2_6_41, w_stg_2_1_42, w_stg_2_7_41, w_stg_2_2_42, w_stg_2_8_41, w_stg_2_3_42, w_stg_2_9_41, w_stg_2_4_42, w_stg_2_10_41, w_stg_2_5_42, w_stg_2_0_43, w_stg_2_6_42, w_stg_2_1_43, w_stg_2_7_42, w_stg_2_2_43, w_stg_2_8_42, w_stg_2_3_43, w_stg_2_9_42, w_stg_2_4_43, w_stg_2_10_42, w_stg_2_5_43, w_stg_2_0_44, w_stg_2_6_43, w_stg_2_1_44, w_stg_2_7_43, w_stg_2_2_44, w_stg_2_8_43, w_stg_2_3_44, w_stg_2_9_43, w_stg_2_4_44, w_stg_2_5_44, w_stg_2_0_45, w_stg_2_6_44, w_stg_2_1_45, w_stg_2_7_44, w_stg_2_2_45, w_stg_2_8_44, w_stg_2_3_45, w_stg_2_9_44, w_stg_2_4_45, w_stg_2_5_45, w_stg_2_0_46, w_stg_2_6_45, w_stg_2_1_46, w_stg_2_7_45, w_stg_2_2_46, w_stg_2_8_45, w_stg_2_3_46, w_stg_2_9_45, w_stg_2_4_46, w_stg_2_5_46, w_stg_2_0_47, w_stg_2_6_46, w_stg_2_1_47, w_stg_2_7_46, w_stg_2_2_47, w_stg_2_8_46, w_stg_2_3_47, w_stg_2_4_47, w_stg_2_0_48, w_stg_2_5_47, w_stg_2_1_48, w_stg_2_6_47, w_stg_2_2_48, w_stg_2_7_47, w_stg_2_3_48, w_stg_2_4_48, w_stg_2_0_49, w_stg_2_5_48, w_stg_2_1_49, w_stg_2_6_48, w_stg_2_2_49, w_stg_2_7_48, w_stg_2_3_49, w_stg_2_4_49, w_stg_2_0_50, w_stg_2_5_49, w_stg_2_1_50, w_stg_2_6_49, w_stg_2_2_50, w_stg_2_7_49, w_stg_2_3_50, w_stg_2_0_51, w_stg_2_4_50, w_stg_2_1_51, w_stg_2_5_50, w_stg_2_2_51, w_stg_2_6_50, w_stg_2_3_51, w_stg_2_0_52, w_stg_2_4_51, w_stg_2_1_52, w_stg_2_5_51, w_stg_2_2_52, w_stg_2_6_51, w_stg_2_3_52, w_stg_2_0_53, w_stg_2_4_52, w_stg_2_1_53, w_stg_2_5_52, w_stg_2_2_53, w_stg_2_3_53, w_stg_2_0_54, w_stg_2_4_53, w_stg_2_1_54, w_stg_2_5_53, w_stg_2_2_54, w_stg_2_3_54, w_stg_2_0_55, w_stg_2_4_54, w_stg_2_1_55, w_stg_2_5_54, w_stg_2_2_55, w_stg_2_3_55, w_stg_2_0_56, w_stg_2_4_55, w_stg_2_1_56, w_stg_2_2_56, w_stg_2_0_57, w_stg_2_3_56, w_stg_2_1_57, w_stg_2_2_57, w_stg_2_0_58, w_stg_2_3_57, w_stg_2_1_58, w_stg_2_2_58, w_stg_2_0_59, w_stg_2_3_58, w_stg_2_1_59, w_stg_2_0_60, w_stg_2_2_59, w_stg_2_1_60, w_stg_2_0_61, w_stg_2_2_60, w_stg_2_1_61, w_stg_2_0_62, w_stg_2_1_62, w_stg_2_0_63;
	wire w_stg_3_0_0, w_stg_3_0_1, w_stg_3_0_2, w_stg_3_0_3, w_stg_3_0_4, w_stg_3_1_4, w_stg_3_0_5, w_stg_3_1_5, w_stg_3_0_6, w_stg_3_1_6, w_stg_3_0_7, w_stg_3_1_7, w_stg_3_0_8, w_stg_3_2_7, w_stg_3_1_8, w_stg_3_0_9, w_stg_3_2_8, w_stg_3_1_9, w_stg_3_0_10, w_stg_3_2_9, w_stg_3_1_10, w_stg_3_2_10, w_stg_3_0_11, w_stg_3_3_10, w_stg_3_1_11, w_stg_3_2_11, w_stg_3_0_12, w_stg_3_3_11, w_stg_3_1_12, w_stg_3_2_12, w_stg_3_0_13, w_stg_3_3_12, w_stg_3_1_13, w_stg_3_2_13, w_stg_3_0_14, w_stg_3_3_13, w_stg_3_1_14, w_stg_3_2_14, w_stg_3_0_15, w_stg_3_3_14, w_stg_3_1_15, w_stg_3_4_14, w_stg_3_2_15, w_stg_3_0_16, w_stg_3_3_15, w_stg_3_1_16, w_stg_3_4_15, w_stg_3_2_16, w_stg_3_0_17, w_stg_3_3_16, w_stg_3_1_17, w_stg_3_4_16, w_stg_3_2_17, w_stg_3_3_17, w_stg_3_0_18, w_stg_3_4_17, w_stg_3_1_18, w_stg_3_5_17, w_stg_3_2_18, w_stg_3_3_18, w_stg_3_0_19, w_stg_3_4_18, w_stg_3_1_19, w_stg_3_5_18, w_stg_3_2_19, w_stg_3_3_19, w_stg_3_0_20, w_stg_3_4_19, w_stg_3_1_20, w_stg_3_5_19, w_stg_3_2_20, w_stg_3_3_20, w_stg_3_0_21, w_stg_3_4_20, w_stg_3_1_21, w_stg_3_5_20, w_stg_3_2_21, w_stg_3_3_21, w_stg_3_0_22, w_stg_3_4_21, w_stg_3_1_22, w_stg_3_5_21, w_stg_3_2_22, w_stg_3_6_21, w_stg_3_3_22, w_stg_3_0_23, w_stg_3_4_22, w_stg_3_1_23, w_stg_3_5_22, w_stg_3_2_23, w_stg_3_6_22, w_stg_3_3_23, w_stg_3_0_24, w_stg_3_4_23, w_stg_3_1_24, w_stg_3_5_23, w_stg_3_2_24, w_stg_3_6_23, w_stg_3_3_24, w_stg_3_4_24, w_stg_3_0_25, w_stg_3_5_24, w_stg_3_1_25, w_stg_3_6_24, w_stg_3_2_25, w_stg_3_7_24, w_stg_3_3_25, w_stg_3_4_25, w_stg_3_0_26, w_stg_3_5_25, w_stg_3_1_26, w_stg_3_6_25, w_stg_3_2_26, w_stg_3_7_25, w_stg_3_3_26, w_stg_3_4_26, w_stg_3_0_27, w_stg_3_5_26, w_stg_3_1_27, w_stg_3_6_26, w_stg_3_2_27, w_stg_3_7_26, w_stg_3_3_27, w_stg_3_4_27, w_stg_3_0_28, w_stg_3_5_27, w_stg_3_1_28, w_stg_3_6_27, w_stg_3_2_28, w_stg_3_7_27, w_stg_3_3_28, w_stg_3_8_27, w_stg_3_4_28, w_stg_3_0_29, w_stg_3_5_28, w_stg_3_1_29, w_stg_3_6_28, w_stg_3_2_29, w_stg_3_7_28, w_stg_3_3_29, w_stg_3_8_28, w_stg_3_4_29, w_stg_3_0_30, w_stg_3_5_29, w_stg_3_1_30, w_stg_3_6_29, w_stg_3_2_30, w_stg_3_7_29, w_stg_3_3_30, w_stg_3_8_29, w_stg_3_4_30, w_stg_3_0_31, w_stg_3_5_30, w_stg_3_1_31, w_stg_3_6_30, w_stg_3_2_31, w_stg_3_7_30, w_stg_3_3_31, w_stg_3_8_30, w_stg_3_4_31, w_stg_3_5_31, w_stg_3_0_32, w_stg_3_6_31, w_stg_3_1_32, w_stg_3_7_31, w_stg_3_2_32, w_stg_3_8_31, w_stg_3_3_32, w_stg_3_9_31, w_stg_3_4_32, w_stg_3_5_32, w_stg_3_0_33, w_stg_3_6_32, w_stg_3_1_33, w_stg_3_7_32, w_stg_3_2_33, w_stg_3_8_32, w_stg_3_3_33, w_stg_3_9_32, w_stg_3_4_33, w_stg_3_5_33, w_stg_3_0_34, w_stg_3_6_33, w_stg_3_1_34, w_stg_3_7_33, w_stg_3_2_34, w_stg_3_8_33, w_stg_3_3_34, w_stg_3_9_33, w_stg_3_4_34, w_stg_3_5_34, w_stg_3_0_35, w_stg_3_6_34, w_stg_3_1_35, w_stg_3_7_34, w_stg_3_2_35, w_stg_3_8_34, w_stg_3_3_35, w_stg_3_9_34, w_stg_3_4_35, w_stg_3_5_35, w_stg_3_0_36, w_stg_3_6_35, w_stg_3_1_36, w_stg_3_7_35, w_stg_3_2_36, w_stg_3_8_35, w_stg_3_3_36, w_stg_3_9_35, w_stg_3_4_36, w_stg_3_5_36, w_stg_3_0_37, w_stg_3_6_36, w_stg_3_1_37, w_stg_3_7_36, w_stg_3_2_37, w_stg_3_8_36, w_stg_3_3_37, w_stg_3_9_36, w_stg_3_4_37, w_stg_3_5_37, w_stg_3_0_38, w_stg_3_6_37, w_stg_3_1_38, w_stg_3_7_37, w_stg_3_2_38, w_stg_3_8_37, w_stg_3_3_38, w_stg_3_9_37, w_stg_3_4_38, w_stg_3_0_39, w_stg_3_5_38, w_stg_3_1_39, w_stg_3_6_38, w_stg_3_2_39, w_stg_3_7_38, w_stg_3_3_39, w_stg_3_4_39, w_stg_3_0_40, w_stg_3_5_39, w_stg_3_1_40, w_stg_3_6_39, w_stg_3_2_40, w_stg_3_7_39, w_stg_3_3_40, w_stg_3_4_40, w_stg_3_0_41, w_stg_3_5_40, w_stg_3_1_41, w_stg_3_6_40, w_stg_3_2_41, w_stg_3_7_40, w_stg_3_3_41, w_stg_3_4_41, w_stg_3_0_42, w_stg_3_5_41, w_stg_3_1_42, w_stg_3_6_41, w_stg_3_2_42, w_stg_3_7_41, w_stg_3_3_42, w_stg_3_4_42, w_stg_3_0_43, w_stg_3_5_42, w_stg_3_1_43, w_stg_3_6_42, w_stg_3_2_43, w_stg_3_7_42, w_stg_3_3_43, w_stg_3_4_43, w_stg_3_0_44, w_stg_3_5_43, w_stg_3_1_44, w_stg_3_6_43, w_stg_3_2_44, w_stg_3_7_43, w_stg_3_3_44, w_stg_3_0_45, w_stg_3_4_44, w_stg_3_1_45, w_stg_3_5_44, w_stg_3_2_45, w_stg_3_6_44, w_stg_3_3_45, w_stg_3_0_46, w_stg_3_4_45, w_stg_3_1_46, w_stg_3_5_45, w_stg_3_2_46, w_stg_3_6_45, w_stg_3_3_46, w_stg_3_0_47, w_stg_3_4_46, w_stg_3_1_47, w_stg_3_5_46, w_stg_3_2_47, w_stg_3_3_47, w_stg_3_0_48, w_stg_3_4_47, w_stg_3_1_48, w_stg_3_5_47, w_stg_3_2_48, w_stg_3_3_48, w_stg_3_0_49, w_stg_3_4_48, w_stg_3_1_49, w_stg_3_5_48, w_stg_3_2_49, w_stg_3_3_49, w_stg_3_0_50, w_stg_3_4_49, w_stg_3_1_50, w_stg_3_5_49, w_stg_3_2_50, w_stg_3_3_50, w_stg_3_0_51, w_stg_3_4_50, w_stg_3_1_51, w_stg_3_5_50, w_stg_3_2_51, w_stg_3_0_52, w_stg_3_3_51, w_stg_3_1_52, w_stg_3_4_51, w_stg_3_2_52, w_stg_3_0_53, w_stg_3_3_52, w_stg_3_1_53, w_stg_3_2_53, w_stg_3_0_54, w_stg_3_3_53, w_stg_3_1_54, w_stg_3_2_54, w_stg_3_0_55, w_stg_3_3_54, w_stg_3_1_55, w_stg_3_2_55, w_stg_3_0_56, w_stg_3_3_55, w_stg_3_1_56, w_stg_3_2_56, w_stg_3_0_57, w_stg_3_3_56, w_stg_3_1_57, w_stg_3_0_58, w_stg_3_2_57, w_stg_3_1_58, w_stg_3_0_59, w_stg_3_2_58, w_stg_3_1_59, w_stg_3_0_60, w_stg_3_1_60, w_stg_3_0_61, w_stg_3_1_61, w_stg_3_0_62, w_stg_3_1_62, w_stg_3_0_63, w_stg_3_1_63;
	wire w_stg_4_0_0, w_stg_4_0_1, w_stg_4_0_2, w_stg_4_0_3, w_stg_4_0_4, w_stg_4_0_5, w_stg_4_1_5, w_stg_4_0_6, w_stg_4_1_6, w_stg_4_0_7, w_stg_4_1_7, w_stg_4_0_8, w_stg_4_1_8, w_stg_4_0_9, w_stg_4_1_9, w_stg_4_0_10, w_stg_4_1_10, w_stg_4_0_11, w_stg_4_2_10, w_stg_4_1_11, w_stg_4_0_12, w_stg_4_2_11, w_stg_4_1_12, w_stg_4_0_13, w_stg_4_2_12, w_stg_4_1_13, w_stg_4_0_14, w_stg_4_2_13, w_stg_4_1_14, w_stg_4_0_15, w_stg_4_2_14, w_stg_4_1_15, w_stg_4_2_15, w_stg_4_0_16, w_stg_4_3_15, w_stg_4_1_16, w_stg_4_2_16, w_stg_4_0_17, w_stg_4_3_16, w_stg_4_1_17, w_stg_4_2_17, w_stg_4_0_18, w_stg_4_3_17, w_stg_4_1_18, w_stg_4_2_18, w_stg_4_0_19, w_stg_4_3_18, w_stg_4_1_19, w_stg_4_2_19, w_stg_4_0_20, w_stg_4_3_19, w_stg_4_1_20, w_stg_4_2_20, w_stg_4_0_21, w_stg_4_3_20, w_stg_4_1_21, w_stg_4_2_21, w_stg_4_0_22, w_stg_4_3_21, w_stg_4_1_22, w_stg_4_4_21, w_stg_4_2_22, w_stg_4_0_23, w_stg_4_3_22, w_stg_4_1_23, w_stg_4_4_22, w_stg_4_2_23, w_stg_4_0_24, w_stg_4_3_23, w_stg_4_1_24, w_stg_4_4_23, w_stg_4_2_24, w_stg_4_0_25, w_stg_4_3_24, w_stg_4_1_25, w_stg_4_4_24, w_stg_4_2_25, w_stg_4_3_25, w_stg_4_0_26, w_stg_4_4_25, w_stg_4_1_26, w_stg_4_5_25, w_stg_4_2_26, w_stg_4_3_26, w_stg_4_0_27, w_stg_4_4_26, w_stg_4_1_27, w_stg_4_5_26, w_stg_4_2_27, w_stg_4_3_27, w_stg_4_0_28, w_stg_4_4_27, w_stg_4_1_28, w_stg_4_5_27, w_stg_4_2_28, w_stg_4_3_28, w_stg_4_0_29, w_stg_4_4_28, w_stg_4_1_29, w_stg_4_5_28, w_stg_4_2_29, w_stg_4_3_29, w_stg_4_0_30, w_stg_4_4_29, w_stg_4_1_30, w_stg_4_5_29, w_stg_4_2_30, w_stg_4_3_30, w_stg_4_0_31, w_stg_4_4_30, w_stg_4_1_31, w_stg_4_5_30, w_stg_4_2_31, w_stg_4_3_31, w_stg_4_0_32, w_stg_4_4_31, w_stg_4_1_32, w_stg_4_5_31, w_stg_4_2_32, w_stg_4_6_31, w_stg_4_3_32, w_stg_4_0_33, w_stg_4_4_32, w_stg_4_1_33, w_stg_4_5_32, w_stg_4_2_33, w_stg_4_6_32, w_stg_4_3_33, w_stg_4_0_34, w_stg_4_4_33, w_stg_4_1_34, w_stg_4_5_33, w_stg_4_2_34, w_stg_4_6_33, w_stg_4_3_34, w_stg_4_0_35, w_stg_4_4_34, w_stg_4_1_35, w_stg_4_5_34, w_stg_4_2_35, w_stg_4_6_34, w_stg_4_3_35, w_stg_4_0_36, w_stg_4_4_35, w_stg_4_1_36, w_stg_4_5_35, w_stg_4_2_36, w_stg_4_6_35, w_stg_4_3_36, w_stg_4_0_37, w_stg_4_4_36, w_stg_4_1_37, w_stg_4_5_36, w_stg_4_2_37, w_stg_4_6_36, w_stg_4_3_37, w_stg_4_0_38, w_stg_4_4_37, w_stg_4_1_38, w_stg_4_5_37, w_stg_4_2_38, w_stg_4_6_37, w_stg_4_3_38, w_stg_4_0_39, w_stg_4_4_38, w_stg_4_1_39, w_stg_4_5_38, w_stg_4_2_39, w_stg_4_3_39, w_stg_4_0_40, w_stg_4_4_39, w_stg_4_1_40, w_stg_4_5_39, w_stg_4_2_40, w_stg_4_3_40, w_stg_4_0_41, w_stg_4_4_40, w_stg_4_1_41, w_stg_4_5_40, w_stg_4_2_41, w_stg_4_3_41, w_stg_4_0_42, w_stg_4_4_41, w_stg_4_1_42, w_stg_4_5_41, w_stg_4_2_42, w_stg_4_3_42, w_stg_4_0_43, w_stg_4_4_42, w_stg_4_1_43, w_stg_4_5_42, w_stg_4_2_43, w_stg_4_3_43, w_stg_4_0_44, w_stg_4_4_43, w_stg_4_1_44, w_stg_4_5_43, w_stg_4_2_44, w_stg_4_3_44, w_stg_4_0_45, w_stg_4_4_44, w_stg_4_1_45, w_stg_4_5_44, w_stg_4_2_45, w_stg_4_0_46, w_stg_4_3_45, w_stg_4_1_46, w_stg_4_4_45, w_stg_4_2_46, w_stg_4_0_47, w_stg_4_3_46, w_stg_4_1_47, w_stg_4_2_47, w_stg_4_0_48, w_stg_4_3_47, w_stg_4_1_48, w_stg_4_2_48, w_stg_4_0_49, w_stg_4_3_48, w_stg_4_1_49, w_stg_4_2_49, w_stg_4_0_50, w_stg_4_3_49, w_stg_4_1_50, w_stg_4_2_50, w_stg_4_0_51, w_stg_4_3_50, w_stg_4_1_51, w_stg_4_2_51, w_stg_4_0_52, w_stg_4_3_51, w_stg_4_1_52, w_stg_4_2_52, w_stg_4_0_53, w_stg_4_3_52, w_stg_4_1_53, w_stg_4_0_54, w_stg_4_2_53, w_stg_4_1_54, w_stg_4_0_55, w_stg_4_2_54, w_stg_4_1_55, w_stg_4_0_56, w_stg_4_2_55, w_stg_4_1_56, w_stg_4_0_57, w_stg_4_2_56, w_stg_4_1_57, w_stg_4_0_58, w_stg_4_1_58, w_stg_4_0_59, w_stg_4_1_59, w_stg_4_0_60, w_stg_4_1_60, w_stg_4_0_61, w_stg_4_1_61, w_stg_4_0_62, w_stg_4_1_62, w_stg_4_0_63, w_stg_4_1_63, w_stg_4_0_64;
	wire w_stg_5_0_0, w_stg_5_0_1, w_stg_5_0_2, w_stg_5_0_3, w_stg_5_0_4, w_stg_5_0_5, w_stg_5_0_6, w_stg_5_1_6, w_stg_5_0_7, w_stg_5_1_7, w_stg_5_0_8, w_stg_5_1_8, w_stg_5_0_9, w_stg_5_1_9, w_stg_5_0_10, w_stg_5_1_10, w_stg_5_0_11, w_stg_5_1_11, w_stg_5_0_12, w_stg_5_1_12, w_stg_5_0_13, w_stg_5_1_13, w_stg_5_0_14, w_stg_5_1_14, w_stg_5_0_15, w_stg_5_1_15, w_stg_5_0_16, w_stg_5_2_15, w_stg_5_1_16, w_stg_5_0_17, w_stg_5_2_16, w_stg_5_1_17, w_stg_5_0_18, w_stg_5_2_17, w_stg_5_1_18, w_stg_5_0_19, w_stg_5_2_18, w_stg_5_1_19, w_stg_5_0_20, w_stg_5_2_19, w_stg_5_1_20, w_stg_5_0_21, w_stg_5_2_20, w_stg_5_1_21, w_stg_5_0_22, w_stg_5_2_21, w_stg_5_1_22, w_stg_5_2_22, w_stg_5_0_23, w_stg_5_3_22, w_stg_5_1_23, w_stg_5_2_23, w_stg_5_0_24, w_stg_5_3_23, w_stg_5_1_24, w_stg_5_2_24, w_stg_5_0_25, w_stg_5_3_24, w_stg_5_1_25, w_stg_5_2_25, w_stg_5_0_26, w_stg_5_3_25, w_stg_5_1_26, w_stg_5_2_26, w_stg_5_0_27, w_stg_5_3_26, w_stg_5_1_27, w_stg_5_2_27, w_stg_5_0_28, w_stg_5_3_27, w_stg_5_1_28, w_stg_5_2_28, w_stg_5_0_29, w_stg_5_3_28, w_stg_5_1_29, w_stg_5_2_29, w_stg_5_0_30, w_stg_5_3_29, w_stg_5_1_30, w_stg_5_2_30, w_stg_5_0_31, w_stg_5_3_30, w_stg_5_1_31, w_stg_5_2_31, w_stg_5_0_32, w_stg_5_3_31, w_stg_5_1_32, w_stg_5_4_31, w_stg_5_2_32, w_stg_5_0_33, w_stg_5_3_32, w_stg_5_1_33, w_stg_5_4_32, w_stg_5_2_33, w_stg_5_0_34, w_stg_5_3_33, w_stg_5_1_34, w_stg_5_4_33, w_stg_5_2_34, w_stg_5_0_35, w_stg_5_3_34, w_stg_5_1_35, w_stg_5_4_34, w_stg_5_2_35, w_stg_5_0_36, w_stg_5_3_35, w_stg_5_1_36, w_stg_5_4_35, w_stg_5_2_36, w_stg_5_0_37, w_stg_5_3_36, w_stg_5_1_37, w_stg_5_4_36, w_stg_5_2_37, w_stg_5_0_38, w_stg_5_3_37, w_stg_5_1_38, w_stg_5_4_37, w_stg_5_2_38, w_stg_5_0_39, w_stg_5_3_38, w_stg_5_1_39, w_stg_5_2_39, w_stg_5_0_40, w_stg_5_3_39, w_stg_5_1_40, w_stg_5_2_40, w_stg_5_0_41, w_stg_5_3_40, w_stg_5_1_41, w_stg_5_2_41, w_stg_5_0_42, w_stg_5_3_41, w_stg_5_1_42, w_stg_5_2_42, w_stg_5_0_43, w_stg_5_3_42, w_stg_5_1_43, w_stg_5_2_43, w_stg_5_0_44, w_stg_5_3_43, w_stg_5_1_44, w_stg_5_2_44, w_stg_5_0_45, w_stg_5_3_44, w_stg_5_1_45, w_stg_5_2_45, w_stg_5_0_46, w_stg_5_3_45, w_stg_5_1_46, w_stg_5_2_46, w_stg_5_0_47, w_stg_5_3_46, w_stg_5_1_47, w_stg_5_0_48, w_stg_5_2_47, w_stg_5_1_48, w_stg_5_0_49, w_stg_5_2_48, w_stg_5_1_49, w_stg_5_0_50, w_stg_5_2_49, w_stg_5_1_50, w_stg_5_0_51, w_stg_5_2_50, w_stg_5_1_51, w_stg_5_0_52, w_stg_5_2_51, w_stg_5_1_52, w_stg_5_0_53, w_stg_5_2_52, w_stg_5_1_53, w_stg_5_0_54, w_stg_5_1_54, w_stg_5_0_55, w_stg_5_1_55, w_stg_5_0_56, w_stg_5_1_56, w_stg_5_0_57, w_stg_5_1_57, w_stg_5_0_58, w_stg_5_1_58, w_stg_5_0_59, w_stg_5_1_59, w_stg_5_0_60, w_stg_5_1_60, w_stg_5_0_61, w_stg_5_1_61, w_stg_5_0_62, w_stg_5_1_62, w_stg_5_0_63, w_stg_5_1_63, w_stg_5_0_64, w_stg_5_1_64;
	wire w_stg_6_0_0, w_stg_6_0_1, w_stg_6_0_2, w_stg_6_0_3, w_stg_6_0_4, w_stg_6_0_5, w_stg_6_0_6, w_stg_6_0_7, w_stg_6_1_7, w_stg_6_0_8, w_stg_6_1_8, w_stg_6_0_9, w_stg_6_1_9, w_stg_6_0_10, w_stg_6_1_10, w_stg_6_0_11, w_stg_6_1_11, w_stg_6_0_12, w_stg_6_1_12, w_stg_6_0_13, w_stg_6_1_13, w_stg_6_0_14, w_stg_6_1_14, w_stg_6_0_15, w_stg_6_1_15, w_stg_6_0_16, w_stg_6_1_16, w_stg_6_0_17, w_stg_6_1_17, w_stg_6_0_18, w_stg_6_1_18, w_stg_6_0_19, w_stg_6_1_19, w_stg_6_0_20, w_stg_6_1_20, w_stg_6_0_21, w_stg_6_1_21, w_stg_6_0_22, w_stg_6_1_22, w_stg_6_0_23, w_stg_6_2_22, w_stg_6_1_23, w_stg_6_0_24, w_stg_6_2_23, w_stg_6_1_24, w_stg_6_0_25, w_stg_6_2_24, w_stg_6_1_25, w_stg_6_0_26, w_stg_6_2_25, w_stg_6_1_26, w_stg_6_0_27, w_stg_6_2_26, w_stg_6_1_27, w_stg_6_0_28, w_stg_6_2_27, w_stg_6_1_28, w_stg_6_0_29, w_stg_6_2_28, w_stg_6_1_29, w_stg_6_0_30, w_stg_6_2_29, w_stg_6_1_30, w_stg_6_0_31, w_stg_6_2_30, w_stg_6_1_31, w_stg_6_0_32, w_stg_6_2_31, w_stg_6_1_32, w_stg_6_2_32, w_stg_6_0_33, w_stg_6_3_32, w_stg_6_1_33, w_stg_6_2_33, w_stg_6_0_34, w_stg_6_3_33, w_stg_6_1_34, w_stg_6_2_34, w_stg_6_0_35, w_stg_6_3_34, w_stg_6_1_35, w_stg_6_2_35, w_stg_6_0_36, w_stg_6_3_35, w_stg_6_1_36, w_stg_6_2_36, w_stg_6_0_37, w_stg_6_3_36, w_stg_6_1_37, w_stg_6_2_37, w_stg_6_0_38, w_stg_6_3_37, w_stg_6_1_38, w_stg_6_2_38, w_stg_6_0_39, w_stg_6_3_38, w_stg_6_1_39, w_stg_6_0_40, w_stg_6_2_39, w_stg_6_1_40, w_stg_6_0_41, w_stg_6_2_40, w_stg_6_1_41, w_stg_6_0_42, w_stg_6_2_41, w_stg_6_1_42, w_stg_6_0_43, w_stg_6_2_42, w_stg_6_1_43, w_stg_6_0_44, w_stg_6_2_43, w_stg_6_1_44, w_stg_6_0_45, w_stg_6_2_44, w_stg_6_1_45, w_stg_6_0_46, w_stg_6_2_45, w_stg_6_1_46, w_stg_6_0_47, w_stg_6_2_46, w_stg_6_1_47, w_stg_6_0_48, w_stg_6_1_48, w_stg_6_0_49, w_stg_6_1_49, w_stg_6_0_50, w_stg_6_1_50, w_stg_6_0_51, w_stg_6_1_51, w_stg_6_0_52, w_stg_6_1_52, w_stg_6_0_53, w_stg_6_1_53, w_stg_6_0_54, w_stg_6_1_54, w_stg_6_0_55, w_stg_6_1_55, w_stg_6_0_56, w_stg_6_1_56, w_stg_6_0_57, w_stg_6_1_57, w_stg_6_0_58, w_stg_6_1_58, w_stg_6_0_59, w_stg_6_1_59, w_stg_6_0_60, w_stg_6_1_60, w_stg_6_0_61, w_stg_6_1_61, w_stg_6_0_62, w_stg_6_1_62, w_stg_6_0_63, w_stg_6_1_63, w_stg_6_0_64, w_stg_6_1_64, w_stg_6_0_65;
	wire w_stg_7_0_0, w_stg_7_0_1, w_stg_7_0_2, w_stg_7_0_3, w_stg_7_0_4, w_stg_7_0_5, w_stg_7_0_6, w_stg_7_0_7, w_stg_7_0_8, w_stg_7_1_8, w_stg_7_0_9, w_stg_7_1_9, w_stg_7_0_10, w_stg_7_1_10, w_stg_7_0_11, w_stg_7_1_11, w_stg_7_0_12, w_stg_7_1_12, w_stg_7_0_13, w_stg_7_1_13, w_stg_7_0_14, w_stg_7_1_14, w_stg_7_0_15, w_stg_7_1_15, w_stg_7_0_16, w_stg_7_1_16, w_stg_7_0_17, w_stg_7_1_17, w_stg_7_0_18, w_stg_7_1_18, w_stg_7_0_19, w_stg_7_1_19, w_stg_7_0_20, w_stg_7_1_20, w_stg_7_0_21, w_stg_7_1_21, w_stg_7_0_22, w_stg_7_1_22, w_stg_7_0_23, w_stg_7_1_23, w_stg_7_0_24, w_stg_7_1_24, w_stg_7_0_25, w_stg_7_1_25, w_stg_7_0_26, w_stg_7_1_26, w_stg_7_0_27, w_stg_7_1_27, w_stg_7_0_28, w_stg_7_1_28, w_stg_7_0_29, w_stg_7_1_29, w_stg_7_0_30, w_stg_7_1_30, w_stg_7_0_31, w_stg_7_1_31, w_stg_7_0_32, w_stg_7_1_32, w_stg_7_0_33, w_stg_7_2_32, w_stg_7_1_33, w_stg_7_0_34, w_stg_7_2_33, w_stg_7_1_34, w_stg_7_0_35, w_stg_7_2_34, w_stg_7_1_35, w_stg_7_0_36, w_stg_7_2_35, w_stg_7_1_36, w_stg_7_0_37, w_stg_7_2_36, w_stg_7_1_37, w_stg_7_0_38, w_stg_7_2_37, w_stg_7_1_38, w_stg_7_0_39, w_stg_7_2_38, w_stg_7_1_39, w_stg_7_0_40, w_stg_7_1_40, w_stg_7_0_41, w_stg_7_1_41, w_stg_7_0_42, w_stg_7_1_42, w_stg_7_0_43, w_stg_7_1_43, w_stg_7_0_44, w_stg_7_1_44, w_stg_7_0_45, w_stg_7_1_45, w_stg_7_0_46, w_stg_7_1_46, w_stg_7_0_47, w_stg_7_1_47, w_stg_7_0_48, w_stg_7_1_48, w_stg_7_0_49, w_stg_7_1_49, w_stg_7_0_50, w_stg_7_1_50, w_stg_7_0_51, w_stg_7_1_51, w_stg_7_0_52, w_stg_7_1_52, w_stg_7_0_53, w_stg_7_1_53, w_stg_7_0_54, w_stg_7_1_54, w_stg_7_0_55, w_stg_7_1_55, w_stg_7_0_56, w_stg_7_1_56, w_stg_7_0_57, w_stg_7_1_57, w_stg_7_0_58, w_stg_7_1_58, w_stg_7_0_59, w_stg_7_1_59, w_stg_7_0_60, w_stg_7_1_60, w_stg_7_0_61, w_stg_7_1_61, w_stg_7_0_62, w_stg_7_1_62, w_stg_7_0_63, w_stg_7_1_63, w_stg_7_0_64, w_stg_7_1_64, w_stg_7_0_65, w_stg_7_1_65;
	wire w_stg_8_0_0, w_stg_8_0_1, w_stg_8_0_2, w_stg_8_0_3, w_stg_8_0_4, w_stg_8_0_5, w_stg_8_0_6, w_stg_8_0_7, w_stg_8_0_8, w_stg_8_0_9, w_stg_8_1_9, w_stg_8_0_10, w_stg_8_1_10, w_stg_8_0_11, w_stg_8_1_11, w_stg_8_0_12, w_stg_8_1_12, w_stg_8_0_13, w_stg_8_1_13, w_stg_8_0_14, w_stg_8_1_14, w_stg_8_0_15, w_stg_8_1_15, w_stg_8_0_16, w_stg_8_1_16, w_stg_8_0_17, w_stg_8_1_17, w_stg_8_0_18, w_stg_8_1_18, w_stg_8_0_19, w_stg_8_1_19, w_stg_8_0_20, w_stg_8_1_20, w_stg_8_0_21, w_stg_8_1_21, w_stg_8_0_22, w_stg_8_1_22, w_stg_8_0_23, w_stg_8_1_23, w_stg_8_0_24, w_stg_8_1_24, w_stg_8_0_25, w_stg_8_1_25, w_stg_8_0_26, w_stg_8_1_26, w_stg_8_0_27, w_stg_8_1_27, w_stg_8_0_28, w_stg_8_1_28, w_stg_8_0_29, w_stg_8_1_29, w_stg_8_0_30, w_stg_8_1_30, w_stg_8_0_31, w_stg_8_1_31, w_stg_8_0_32, w_stg_8_1_32, w_stg_8_0_33, w_stg_8_1_33, w_stg_8_0_34, w_stg_8_1_34, w_stg_8_0_35, w_stg_8_1_35, w_stg_8_0_36, w_stg_8_1_36, w_stg_8_0_37, w_stg_8_1_37, w_stg_8_0_38, w_stg_8_1_38, w_stg_8_0_39, w_stg_8_1_39, w_stg_8_0_40, w_stg_8_1_40, w_stg_8_0_41, w_stg_8_1_41, w_stg_8_0_42, w_stg_8_1_42, w_stg_8_0_43, w_stg_8_1_43, w_stg_8_0_44, w_stg_8_1_44, w_stg_8_0_45, w_stg_8_1_45, w_stg_8_0_46, w_stg_8_1_46, w_stg_8_0_47, w_stg_8_1_47, w_stg_8_0_48, w_stg_8_1_48, w_stg_8_0_49, w_stg_8_1_49, w_stg_8_0_50, w_stg_8_1_50, w_stg_8_0_51, w_stg_8_1_51, w_stg_8_0_52, w_stg_8_1_52, w_stg_8_0_53, w_stg_8_1_53, w_stg_8_0_54, w_stg_8_1_54, w_stg_8_0_55, w_stg_8_1_55, w_stg_8_0_56, w_stg_8_1_56, w_stg_8_0_57, w_stg_8_1_57, w_stg_8_0_58, w_stg_8_1_58, w_stg_8_0_59, w_stg_8_1_59, w_stg_8_0_60, w_stg_8_1_60, w_stg_8_0_61, w_stg_8_1_61, w_stg_8_0_62, w_stg_8_1_62, w_stg_8_0_63, w_stg_8_1_63, w_stg_8_0_64, w_stg_8_1_64, w_stg_8_0_65, w_stg_8_1_65, w_stg_8_0_66;


	and stg_0_0_0(w_stg_0_0_0, data_operandA[0], data_operandB[0]);
	and stg_0_0_1(w_stg_0_0_1, data_operandA[1], data_operandB[0]);
	and stg_0_0_2(w_stg_0_0_2, data_operandA[2], data_operandB[0]);
	and stg_0_0_3(w_stg_0_0_3, data_operandA[3], data_operandB[0]);
	and stg_0_0_4(w_stg_0_0_4, data_operandA[4], data_operandB[0]);
	and stg_0_0_5(w_stg_0_0_5, data_operandA[5], data_operandB[0]);
	and stg_0_0_6(w_stg_0_0_6, data_operandA[6], data_operandB[0]);
	and stg_0_0_7(w_stg_0_0_7, data_operandA[7], data_operandB[0]);
	and stg_0_0_8(w_stg_0_0_8, data_operandA[8], data_operandB[0]);
	and stg_0_0_9(w_stg_0_0_9, data_operandA[9], data_operandB[0]);
	and stg_0_0_10(w_stg_0_0_10, data_operandA[10], data_operandB[0]);
	and stg_0_0_11(w_stg_0_0_11, data_operandA[11], data_operandB[0]);
	and stg_0_0_12(w_stg_0_0_12, data_operandA[12], data_operandB[0]);
	and stg_0_0_13(w_stg_0_0_13, data_operandA[13], data_operandB[0]);
	and stg_0_0_14(w_stg_0_0_14, data_operandA[14], data_operandB[0]);
	and stg_0_0_15(w_stg_0_0_15, data_operandA[15], data_operandB[0]);
	and stg_0_0_16(w_stg_0_0_16, data_operandA[16], data_operandB[0]);
	and stg_0_0_17(w_stg_0_0_17, data_operandA[17], data_operandB[0]);
	and stg_0_0_18(w_stg_0_0_18, data_operandA[18], data_operandB[0]);
	and stg_0_0_19(w_stg_0_0_19, data_operandA[19], data_operandB[0]);
	and stg_0_0_20(w_stg_0_0_20, data_operandA[20], data_operandB[0]);
	and stg_0_0_21(w_stg_0_0_21, data_operandA[21], data_operandB[0]);
	and stg_0_0_22(w_stg_0_0_22, data_operandA[22], data_operandB[0]);
	and stg_0_0_23(w_stg_0_0_23, data_operandA[23], data_operandB[0]);
	and stg_0_0_24(w_stg_0_0_24, data_operandA[24], data_operandB[0]);
	and stg_0_0_25(w_stg_0_0_25, data_operandA[25], data_operandB[0]);
	and stg_0_0_26(w_stg_0_0_26, data_operandA[26], data_operandB[0]);
	and stg_0_0_27(w_stg_0_0_27, data_operandA[27], data_operandB[0]);
	and stg_0_0_28(w_stg_0_0_28, data_operandA[28], data_operandB[0]);
	and stg_0_0_29(w_stg_0_0_29, data_operandA[29], data_operandB[0]);
	and stg_0_0_30(w_stg_0_0_30, data_operandA[30], data_operandB[0]);
	and stg_0_0_31(w_stg_0_0_31, data_operandA[31], data_operandB[0]);
	and stg_0_1_1(w_stg_0_1_1, data_operandA[0], data_operandB[1]);
	and stg_0_1_2(w_stg_0_1_2, data_operandA[1], data_operandB[1]);
	and stg_0_1_3(w_stg_0_1_3, data_operandA[2], data_operandB[1]);
	and stg_0_1_4(w_stg_0_1_4, data_operandA[3], data_operandB[1]);
	and stg_0_1_5(w_stg_0_1_5, data_operandA[4], data_operandB[1]);
	and stg_0_1_6(w_stg_0_1_6, data_operandA[5], data_operandB[1]);
	and stg_0_1_7(w_stg_0_1_7, data_operandA[6], data_operandB[1]);
	and stg_0_1_8(w_stg_0_1_8, data_operandA[7], data_operandB[1]);
	and stg_0_1_9(w_stg_0_1_9, data_operandA[8], data_operandB[1]);
	and stg_0_1_10(w_stg_0_1_10, data_operandA[9], data_operandB[1]);
	and stg_0_1_11(w_stg_0_1_11, data_operandA[10], data_operandB[1]);
	and stg_0_1_12(w_stg_0_1_12, data_operandA[11], data_operandB[1]);
	and stg_0_1_13(w_stg_0_1_13, data_operandA[12], data_operandB[1]);
	and stg_0_1_14(w_stg_0_1_14, data_operandA[13], data_operandB[1]);
	and stg_0_1_15(w_stg_0_1_15, data_operandA[14], data_operandB[1]);
	and stg_0_1_16(w_stg_0_1_16, data_operandA[15], data_operandB[1]);
	and stg_0_1_17(w_stg_0_1_17, data_operandA[16], data_operandB[1]);
	and stg_0_1_18(w_stg_0_1_18, data_operandA[17], data_operandB[1]);
	and stg_0_1_19(w_stg_0_1_19, data_operandA[18], data_operandB[1]);
	and stg_0_1_20(w_stg_0_1_20, data_operandA[19], data_operandB[1]);
	and stg_0_1_21(w_stg_0_1_21, data_operandA[20], data_operandB[1]);
	and stg_0_1_22(w_stg_0_1_22, data_operandA[21], data_operandB[1]);
	and stg_0_1_23(w_stg_0_1_23, data_operandA[22], data_operandB[1]);
	and stg_0_1_24(w_stg_0_1_24, data_operandA[23], data_operandB[1]);
	and stg_0_1_25(w_stg_0_1_25, data_operandA[24], data_operandB[1]);
	and stg_0_1_26(w_stg_0_1_26, data_operandA[25], data_operandB[1]);
	and stg_0_1_27(w_stg_0_1_27, data_operandA[26], data_operandB[1]);
	and stg_0_1_28(w_stg_0_1_28, data_operandA[27], data_operandB[1]);
	and stg_0_1_29(w_stg_0_1_29, data_operandA[28], data_operandB[1]);
	and stg_0_1_30(w_stg_0_1_30, data_operandA[29], data_operandB[1]);
	and stg_0_1_31(w_stg_0_1_31, data_operandA[30], data_operandB[1]);
	and stg_0_1_32(w_stg_0_1_32, data_operandA[31], data_operandB[1]);
	and stg_0_2_2(w_stg_0_2_2, data_operandA[0], data_operandB[2]);
	and stg_0_2_3(w_stg_0_2_3, data_operandA[1], data_operandB[2]);
	and stg_0_2_4(w_stg_0_2_4, data_operandA[2], data_operandB[2]);
	and stg_0_2_5(w_stg_0_2_5, data_operandA[3], data_operandB[2]);
	and stg_0_2_6(w_stg_0_2_6, data_operandA[4], data_operandB[2]);
	and stg_0_2_7(w_stg_0_2_7, data_operandA[5], data_operandB[2]);
	and stg_0_2_8(w_stg_0_2_8, data_operandA[6], data_operandB[2]);
	and stg_0_2_9(w_stg_0_2_9, data_operandA[7], data_operandB[2]);
	and stg_0_2_10(w_stg_0_2_10, data_operandA[8], data_operandB[2]);
	and stg_0_2_11(w_stg_0_2_11, data_operandA[9], data_operandB[2]);
	and stg_0_2_12(w_stg_0_2_12, data_operandA[10], data_operandB[2]);
	and stg_0_2_13(w_stg_0_2_13, data_operandA[11], data_operandB[2]);
	and stg_0_2_14(w_stg_0_2_14, data_operandA[12], data_operandB[2]);
	and stg_0_2_15(w_stg_0_2_15, data_operandA[13], data_operandB[2]);
	and stg_0_2_16(w_stg_0_2_16, data_operandA[14], data_operandB[2]);
	and stg_0_2_17(w_stg_0_2_17, data_operandA[15], data_operandB[2]);
	and stg_0_2_18(w_stg_0_2_18, data_operandA[16], data_operandB[2]);
	and stg_0_2_19(w_stg_0_2_19, data_operandA[17], data_operandB[2]);
	and stg_0_2_20(w_stg_0_2_20, data_operandA[18], data_operandB[2]);
	and stg_0_2_21(w_stg_0_2_21, data_operandA[19], data_operandB[2]);
	and stg_0_2_22(w_stg_0_2_22, data_operandA[20], data_operandB[2]);
	and stg_0_2_23(w_stg_0_2_23, data_operandA[21], data_operandB[2]);
	and stg_0_2_24(w_stg_0_2_24, data_operandA[22], data_operandB[2]);
	and stg_0_2_25(w_stg_0_2_25, data_operandA[23], data_operandB[2]);
	and stg_0_2_26(w_stg_0_2_26, data_operandA[24], data_operandB[2]);
	and stg_0_2_27(w_stg_0_2_27, data_operandA[25], data_operandB[2]);
	and stg_0_2_28(w_stg_0_2_28, data_operandA[26], data_operandB[2]);
	and stg_0_2_29(w_stg_0_2_29, data_operandA[27], data_operandB[2]);
	and stg_0_2_30(w_stg_0_2_30, data_operandA[28], data_operandB[2]);
	and stg_0_2_31(w_stg_0_2_31, data_operandA[29], data_operandB[2]);
	and stg_0_2_32(w_stg_0_2_32, data_operandA[30], data_operandB[2]);
	and stg_0_2_33(w_stg_0_2_33, data_operandA[31], data_operandB[2]);
	and stg_0_3_3(w_stg_0_3_3, data_operandA[0], data_operandB[3]);
	and stg_0_3_4(w_stg_0_3_4, data_operandA[1], data_operandB[3]);
	and stg_0_3_5(w_stg_0_3_5, data_operandA[2], data_operandB[3]);
	and stg_0_3_6(w_stg_0_3_6, data_operandA[3], data_operandB[3]);
	and stg_0_3_7(w_stg_0_3_7, data_operandA[4], data_operandB[3]);
	and stg_0_3_8(w_stg_0_3_8, data_operandA[5], data_operandB[3]);
	and stg_0_3_9(w_stg_0_3_9, data_operandA[6], data_operandB[3]);
	and stg_0_3_10(w_stg_0_3_10, data_operandA[7], data_operandB[3]);
	and stg_0_3_11(w_stg_0_3_11, data_operandA[8], data_operandB[3]);
	and stg_0_3_12(w_stg_0_3_12, data_operandA[9], data_operandB[3]);
	and stg_0_3_13(w_stg_0_3_13, data_operandA[10], data_operandB[3]);
	and stg_0_3_14(w_stg_0_3_14, data_operandA[11], data_operandB[3]);
	and stg_0_3_15(w_stg_0_3_15, data_operandA[12], data_operandB[3]);
	and stg_0_3_16(w_stg_0_3_16, data_operandA[13], data_operandB[3]);
	and stg_0_3_17(w_stg_0_3_17, data_operandA[14], data_operandB[3]);
	and stg_0_3_18(w_stg_0_3_18, data_operandA[15], data_operandB[3]);
	and stg_0_3_19(w_stg_0_3_19, data_operandA[16], data_operandB[3]);
	and stg_0_3_20(w_stg_0_3_20, data_operandA[17], data_operandB[3]);
	and stg_0_3_21(w_stg_0_3_21, data_operandA[18], data_operandB[3]);
	and stg_0_3_22(w_stg_0_3_22, data_operandA[19], data_operandB[3]);
	and stg_0_3_23(w_stg_0_3_23, data_operandA[20], data_operandB[3]);
	and stg_0_3_24(w_stg_0_3_24, data_operandA[21], data_operandB[3]);
	and stg_0_3_25(w_stg_0_3_25, data_operandA[22], data_operandB[3]);
	and stg_0_3_26(w_stg_0_3_26, data_operandA[23], data_operandB[3]);
	and stg_0_3_27(w_stg_0_3_27, data_operandA[24], data_operandB[3]);
	and stg_0_3_28(w_stg_0_3_28, data_operandA[25], data_operandB[3]);
	and stg_0_3_29(w_stg_0_3_29, data_operandA[26], data_operandB[3]);
	and stg_0_3_30(w_stg_0_3_30, data_operandA[27], data_operandB[3]);
	and stg_0_3_31(w_stg_0_3_31, data_operandA[28], data_operandB[3]);
	and stg_0_3_32(w_stg_0_3_32, data_operandA[29], data_operandB[3]);
	and stg_0_3_33(w_stg_0_3_33, data_operandA[30], data_operandB[3]);
	and stg_0_3_34(w_stg_0_3_34, data_operandA[31], data_operandB[3]);
	and stg_0_4_4(w_stg_0_4_4, data_operandA[0], data_operandB[4]);
	and stg_0_4_5(w_stg_0_4_5, data_operandA[1], data_operandB[4]);
	and stg_0_4_6(w_stg_0_4_6, data_operandA[2], data_operandB[4]);
	and stg_0_4_7(w_stg_0_4_7, data_operandA[3], data_operandB[4]);
	and stg_0_4_8(w_stg_0_4_8, data_operandA[4], data_operandB[4]);
	and stg_0_4_9(w_stg_0_4_9, data_operandA[5], data_operandB[4]);
	and stg_0_4_10(w_stg_0_4_10, data_operandA[6], data_operandB[4]);
	and stg_0_4_11(w_stg_0_4_11, data_operandA[7], data_operandB[4]);
	and stg_0_4_12(w_stg_0_4_12, data_operandA[8], data_operandB[4]);
	and stg_0_4_13(w_stg_0_4_13, data_operandA[9], data_operandB[4]);
	and stg_0_4_14(w_stg_0_4_14, data_operandA[10], data_operandB[4]);
	and stg_0_4_15(w_stg_0_4_15, data_operandA[11], data_operandB[4]);
	and stg_0_4_16(w_stg_0_4_16, data_operandA[12], data_operandB[4]);
	and stg_0_4_17(w_stg_0_4_17, data_operandA[13], data_operandB[4]);
	and stg_0_4_18(w_stg_0_4_18, data_operandA[14], data_operandB[4]);
	and stg_0_4_19(w_stg_0_4_19, data_operandA[15], data_operandB[4]);
	and stg_0_4_20(w_stg_0_4_20, data_operandA[16], data_operandB[4]);
	and stg_0_4_21(w_stg_0_4_21, data_operandA[17], data_operandB[4]);
	and stg_0_4_22(w_stg_0_4_22, data_operandA[18], data_operandB[4]);
	and stg_0_4_23(w_stg_0_4_23, data_operandA[19], data_operandB[4]);
	and stg_0_4_24(w_stg_0_4_24, data_operandA[20], data_operandB[4]);
	and stg_0_4_25(w_stg_0_4_25, data_operandA[21], data_operandB[4]);
	and stg_0_4_26(w_stg_0_4_26, data_operandA[22], data_operandB[4]);
	and stg_0_4_27(w_stg_0_4_27, data_operandA[23], data_operandB[4]);
	and stg_0_4_28(w_stg_0_4_28, data_operandA[24], data_operandB[4]);
	and stg_0_4_29(w_stg_0_4_29, data_operandA[25], data_operandB[4]);
	and stg_0_4_30(w_stg_0_4_30, data_operandA[26], data_operandB[4]);
	and stg_0_4_31(w_stg_0_4_31, data_operandA[27], data_operandB[4]);
	and stg_0_4_32(w_stg_0_4_32, data_operandA[28], data_operandB[4]);
	and stg_0_4_33(w_stg_0_4_33, data_operandA[29], data_operandB[4]);
	and stg_0_4_34(w_stg_0_4_34, data_operandA[30], data_operandB[4]);
	and stg_0_4_35(w_stg_0_4_35, data_operandA[31], data_operandB[4]);
	and stg_0_5_5(w_stg_0_5_5, data_operandA[0], data_operandB[5]);
	and stg_0_5_6(w_stg_0_5_6, data_operandA[1], data_operandB[5]);
	and stg_0_5_7(w_stg_0_5_7, data_operandA[2], data_operandB[5]);
	and stg_0_5_8(w_stg_0_5_8, data_operandA[3], data_operandB[5]);
	and stg_0_5_9(w_stg_0_5_9, data_operandA[4], data_operandB[5]);
	and stg_0_5_10(w_stg_0_5_10, data_operandA[5], data_operandB[5]);
	and stg_0_5_11(w_stg_0_5_11, data_operandA[6], data_operandB[5]);
	and stg_0_5_12(w_stg_0_5_12, data_operandA[7], data_operandB[5]);
	and stg_0_5_13(w_stg_0_5_13, data_operandA[8], data_operandB[5]);
	and stg_0_5_14(w_stg_0_5_14, data_operandA[9], data_operandB[5]);
	and stg_0_5_15(w_stg_0_5_15, data_operandA[10], data_operandB[5]);
	and stg_0_5_16(w_stg_0_5_16, data_operandA[11], data_operandB[5]);
	and stg_0_5_17(w_stg_0_5_17, data_operandA[12], data_operandB[5]);
	and stg_0_5_18(w_stg_0_5_18, data_operandA[13], data_operandB[5]);
	and stg_0_5_19(w_stg_0_5_19, data_operandA[14], data_operandB[5]);
	and stg_0_5_20(w_stg_0_5_20, data_operandA[15], data_operandB[5]);
	and stg_0_5_21(w_stg_0_5_21, data_operandA[16], data_operandB[5]);
	and stg_0_5_22(w_stg_0_5_22, data_operandA[17], data_operandB[5]);
	and stg_0_5_23(w_stg_0_5_23, data_operandA[18], data_operandB[5]);
	and stg_0_5_24(w_stg_0_5_24, data_operandA[19], data_operandB[5]);
	and stg_0_5_25(w_stg_0_5_25, data_operandA[20], data_operandB[5]);
	and stg_0_5_26(w_stg_0_5_26, data_operandA[21], data_operandB[5]);
	and stg_0_5_27(w_stg_0_5_27, data_operandA[22], data_operandB[5]);
	and stg_0_5_28(w_stg_0_5_28, data_operandA[23], data_operandB[5]);
	and stg_0_5_29(w_stg_0_5_29, data_operandA[24], data_operandB[5]);
	and stg_0_5_30(w_stg_0_5_30, data_operandA[25], data_operandB[5]);
	and stg_0_5_31(w_stg_0_5_31, data_operandA[26], data_operandB[5]);
	and stg_0_5_32(w_stg_0_5_32, data_operandA[27], data_operandB[5]);
	and stg_0_5_33(w_stg_0_5_33, data_operandA[28], data_operandB[5]);
	and stg_0_5_34(w_stg_0_5_34, data_operandA[29], data_operandB[5]);
	and stg_0_5_35(w_stg_0_5_35, data_operandA[30], data_operandB[5]);
	and stg_0_5_36(w_stg_0_5_36, data_operandA[31], data_operandB[5]);
	and stg_0_6_6(w_stg_0_6_6, data_operandA[0], data_operandB[6]);
	and stg_0_6_7(w_stg_0_6_7, data_operandA[1], data_operandB[6]);
	and stg_0_6_8(w_stg_0_6_8, data_operandA[2], data_operandB[6]);
	and stg_0_6_9(w_stg_0_6_9, data_operandA[3], data_operandB[6]);
	and stg_0_6_10(w_stg_0_6_10, data_operandA[4], data_operandB[6]);
	and stg_0_6_11(w_stg_0_6_11, data_operandA[5], data_operandB[6]);
	and stg_0_6_12(w_stg_0_6_12, data_operandA[6], data_operandB[6]);
	and stg_0_6_13(w_stg_0_6_13, data_operandA[7], data_operandB[6]);
	and stg_0_6_14(w_stg_0_6_14, data_operandA[8], data_operandB[6]);
	and stg_0_6_15(w_stg_0_6_15, data_operandA[9], data_operandB[6]);
	and stg_0_6_16(w_stg_0_6_16, data_operandA[10], data_operandB[6]);
	and stg_0_6_17(w_stg_0_6_17, data_operandA[11], data_operandB[6]);
	and stg_0_6_18(w_stg_0_6_18, data_operandA[12], data_operandB[6]);
	and stg_0_6_19(w_stg_0_6_19, data_operandA[13], data_operandB[6]);
	and stg_0_6_20(w_stg_0_6_20, data_operandA[14], data_operandB[6]);
	and stg_0_6_21(w_stg_0_6_21, data_operandA[15], data_operandB[6]);
	and stg_0_6_22(w_stg_0_6_22, data_operandA[16], data_operandB[6]);
	and stg_0_6_23(w_stg_0_6_23, data_operandA[17], data_operandB[6]);
	and stg_0_6_24(w_stg_0_6_24, data_operandA[18], data_operandB[6]);
	and stg_0_6_25(w_stg_0_6_25, data_operandA[19], data_operandB[6]);
	and stg_0_6_26(w_stg_0_6_26, data_operandA[20], data_operandB[6]);
	and stg_0_6_27(w_stg_0_6_27, data_operandA[21], data_operandB[6]);
	and stg_0_6_28(w_stg_0_6_28, data_operandA[22], data_operandB[6]);
	and stg_0_6_29(w_stg_0_6_29, data_operandA[23], data_operandB[6]);
	and stg_0_6_30(w_stg_0_6_30, data_operandA[24], data_operandB[6]);
	and stg_0_6_31(w_stg_0_6_31, data_operandA[25], data_operandB[6]);
	and stg_0_6_32(w_stg_0_6_32, data_operandA[26], data_operandB[6]);
	and stg_0_6_33(w_stg_0_6_33, data_operandA[27], data_operandB[6]);
	and stg_0_6_34(w_stg_0_6_34, data_operandA[28], data_operandB[6]);
	and stg_0_6_35(w_stg_0_6_35, data_operandA[29], data_operandB[6]);
	and stg_0_6_36(w_stg_0_6_36, data_operandA[30], data_operandB[6]);
	and stg_0_6_37(w_stg_0_6_37, data_operandA[31], data_operandB[6]);
	and stg_0_7_7(w_stg_0_7_7, data_operandA[0], data_operandB[7]);
	and stg_0_7_8(w_stg_0_7_8, data_operandA[1], data_operandB[7]);
	and stg_0_7_9(w_stg_0_7_9, data_operandA[2], data_operandB[7]);
	and stg_0_7_10(w_stg_0_7_10, data_operandA[3], data_operandB[7]);
	and stg_0_7_11(w_stg_0_7_11, data_operandA[4], data_operandB[7]);
	and stg_0_7_12(w_stg_0_7_12, data_operandA[5], data_operandB[7]);
	and stg_0_7_13(w_stg_0_7_13, data_operandA[6], data_operandB[7]);
	and stg_0_7_14(w_stg_0_7_14, data_operandA[7], data_operandB[7]);
	and stg_0_7_15(w_stg_0_7_15, data_operandA[8], data_operandB[7]);
	and stg_0_7_16(w_stg_0_7_16, data_operandA[9], data_operandB[7]);
	and stg_0_7_17(w_stg_0_7_17, data_operandA[10], data_operandB[7]);
	and stg_0_7_18(w_stg_0_7_18, data_operandA[11], data_operandB[7]);
	and stg_0_7_19(w_stg_0_7_19, data_operandA[12], data_operandB[7]);
	and stg_0_7_20(w_stg_0_7_20, data_operandA[13], data_operandB[7]);
	and stg_0_7_21(w_stg_0_7_21, data_operandA[14], data_operandB[7]);
	and stg_0_7_22(w_stg_0_7_22, data_operandA[15], data_operandB[7]);
	and stg_0_7_23(w_stg_0_7_23, data_operandA[16], data_operandB[7]);
	and stg_0_7_24(w_stg_0_7_24, data_operandA[17], data_operandB[7]);
	and stg_0_7_25(w_stg_0_7_25, data_operandA[18], data_operandB[7]);
	and stg_0_7_26(w_stg_0_7_26, data_operandA[19], data_operandB[7]);
	and stg_0_7_27(w_stg_0_7_27, data_operandA[20], data_operandB[7]);
	and stg_0_7_28(w_stg_0_7_28, data_operandA[21], data_operandB[7]);
	and stg_0_7_29(w_stg_0_7_29, data_operandA[22], data_operandB[7]);
	and stg_0_7_30(w_stg_0_7_30, data_operandA[23], data_operandB[7]);
	and stg_0_7_31(w_stg_0_7_31, data_operandA[24], data_operandB[7]);
	and stg_0_7_32(w_stg_0_7_32, data_operandA[25], data_operandB[7]);
	and stg_0_7_33(w_stg_0_7_33, data_operandA[26], data_operandB[7]);
	and stg_0_7_34(w_stg_0_7_34, data_operandA[27], data_operandB[7]);
	and stg_0_7_35(w_stg_0_7_35, data_operandA[28], data_operandB[7]);
	and stg_0_7_36(w_stg_0_7_36, data_operandA[29], data_operandB[7]);
	and stg_0_7_37(w_stg_0_7_37, data_operandA[30], data_operandB[7]);
	and stg_0_7_38(w_stg_0_7_38, data_operandA[31], data_operandB[7]);
	and stg_0_8_8(w_stg_0_8_8, data_operandA[0], data_operandB[8]);
	and stg_0_8_9(w_stg_0_8_9, data_operandA[1], data_operandB[8]);
	and stg_0_8_10(w_stg_0_8_10, data_operandA[2], data_operandB[8]);
	and stg_0_8_11(w_stg_0_8_11, data_operandA[3], data_operandB[8]);
	and stg_0_8_12(w_stg_0_8_12, data_operandA[4], data_operandB[8]);
	and stg_0_8_13(w_stg_0_8_13, data_operandA[5], data_operandB[8]);
	and stg_0_8_14(w_stg_0_8_14, data_operandA[6], data_operandB[8]);
	and stg_0_8_15(w_stg_0_8_15, data_operandA[7], data_operandB[8]);
	and stg_0_8_16(w_stg_0_8_16, data_operandA[8], data_operandB[8]);
	and stg_0_8_17(w_stg_0_8_17, data_operandA[9], data_operandB[8]);
	and stg_0_8_18(w_stg_0_8_18, data_operandA[10], data_operandB[8]);
	and stg_0_8_19(w_stg_0_8_19, data_operandA[11], data_operandB[8]);
	and stg_0_8_20(w_stg_0_8_20, data_operandA[12], data_operandB[8]);
	and stg_0_8_21(w_stg_0_8_21, data_operandA[13], data_operandB[8]);
	and stg_0_8_22(w_stg_0_8_22, data_operandA[14], data_operandB[8]);
	and stg_0_8_23(w_stg_0_8_23, data_operandA[15], data_operandB[8]);
	and stg_0_8_24(w_stg_0_8_24, data_operandA[16], data_operandB[8]);
	and stg_0_8_25(w_stg_0_8_25, data_operandA[17], data_operandB[8]);
	and stg_0_8_26(w_stg_0_8_26, data_operandA[18], data_operandB[8]);
	and stg_0_8_27(w_stg_0_8_27, data_operandA[19], data_operandB[8]);
	and stg_0_8_28(w_stg_0_8_28, data_operandA[20], data_operandB[8]);
	and stg_0_8_29(w_stg_0_8_29, data_operandA[21], data_operandB[8]);
	and stg_0_8_30(w_stg_0_8_30, data_operandA[22], data_operandB[8]);
	and stg_0_8_31(w_stg_0_8_31, data_operandA[23], data_operandB[8]);
	and stg_0_8_32(w_stg_0_8_32, data_operandA[24], data_operandB[8]);
	and stg_0_8_33(w_stg_0_8_33, data_operandA[25], data_operandB[8]);
	and stg_0_8_34(w_stg_0_8_34, data_operandA[26], data_operandB[8]);
	and stg_0_8_35(w_stg_0_8_35, data_operandA[27], data_operandB[8]);
	and stg_0_8_36(w_stg_0_8_36, data_operandA[28], data_operandB[8]);
	and stg_0_8_37(w_stg_0_8_37, data_operandA[29], data_operandB[8]);
	and stg_0_8_38(w_stg_0_8_38, data_operandA[30], data_operandB[8]);
	and stg_0_8_39(w_stg_0_8_39, data_operandA[31], data_operandB[8]);
	and stg_0_9_9(w_stg_0_9_9, data_operandA[0], data_operandB[9]);
	and stg_0_9_10(w_stg_0_9_10, data_operandA[1], data_operandB[9]);
	and stg_0_9_11(w_stg_0_9_11, data_operandA[2], data_operandB[9]);
	and stg_0_9_12(w_stg_0_9_12, data_operandA[3], data_operandB[9]);
	and stg_0_9_13(w_stg_0_9_13, data_operandA[4], data_operandB[9]);
	and stg_0_9_14(w_stg_0_9_14, data_operandA[5], data_operandB[9]);
	and stg_0_9_15(w_stg_0_9_15, data_operandA[6], data_operandB[9]);
	and stg_0_9_16(w_stg_0_9_16, data_operandA[7], data_operandB[9]);
	and stg_0_9_17(w_stg_0_9_17, data_operandA[8], data_operandB[9]);
	and stg_0_9_18(w_stg_0_9_18, data_operandA[9], data_operandB[9]);
	and stg_0_9_19(w_stg_0_9_19, data_operandA[10], data_operandB[9]);
	and stg_0_9_20(w_stg_0_9_20, data_operandA[11], data_operandB[9]);
	and stg_0_9_21(w_stg_0_9_21, data_operandA[12], data_operandB[9]);
	and stg_0_9_22(w_stg_0_9_22, data_operandA[13], data_operandB[9]);
	and stg_0_9_23(w_stg_0_9_23, data_operandA[14], data_operandB[9]);
	and stg_0_9_24(w_stg_0_9_24, data_operandA[15], data_operandB[9]);
	and stg_0_9_25(w_stg_0_9_25, data_operandA[16], data_operandB[9]);
	and stg_0_9_26(w_stg_0_9_26, data_operandA[17], data_operandB[9]);
	and stg_0_9_27(w_stg_0_9_27, data_operandA[18], data_operandB[9]);
	and stg_0_9_28(w_stg_0_9_28, data_operandA[19], data_operandB[9]);
	and stg_0_9_29(w_stg_0_9_29, data_operandA[20], data_operandB[9]);
	and stg_0_9_30(w_stg_0_9_30, data_operandA[21], data_operandB[9]);
	and stg_0_9_31(w_stg_0_9_31, data_operandA[22], data_operandB[9]);
	and stg_0_9_32(w_stg_0_9_32, data_operandA[23], data_operandB[9]);
	and stg_0_9_33(w_stg_0_9_33, data_operandA[24], data_operandB[9]);
	and stg_0_9_34(w_stg_0_9_34, data_operandA[25], data_operandB[9]);
	and stg_0_9_35(w_stg_0_9_35, data_operandA[26], data_operandB[9]);
	and stg_0_9_36(w_stg_0_9_36, data_operandA[27], data_operandB[9]);
	and stg_0_9_37(w_stg_0_9_37, data_operandA[28], data_operandB[9]);
	and stg_0_9_38(w_stg_0_9_38, data_operandA[29], data_operandB[9]);
	and stg_0_9_39(w_stg_0_9_39, data_operandA[30], data_operandB[9]);
	and stg_0_9_40(w_stg_0_9_40, data_operandA[31], data_operandB[9]);
	and stg_0_10_10(w_stg_0_10_10, data_operandA[0], data_operandB[10]);
	and stg_0_10_11(w_stg_0_10_11, data_operandA[1], data_operandB[10]);
	and stg_0_10_12(w_stg_0_10_12, data_operandA[2], data_operandB[10]);
	and stg_0_10_13(w_stg_0_10_13, data_operandA[3], data_operandB[10]);
	and stg_0_10_14(w_stg_0_10_14, data_operandA[4], data_operandB[10]);
	and stg_0_10_15(w_stg_0_10_15, data_operandA[5], data_operandB[10]);
	and stg_0_10_16(w_stg_0_10_16, data_operandA[6], data_operandB[10]);
	and stg_0_10_17(w_stg_0_10_17, data_operandA[7], data_operandB[10]);
	and stg_0_10_18(w_stg_0_10_18, data_operandA[8], data_operandB[10]);
	and stg_0_10_19(w_stg_0_10_19, data_operandA[9], data_operandB[10]);
	and stg_0_10_20(w_stg_0_10_20, data_operandA[10], data_operandB[10]);
	and stg_0_10_21(w_stg_0_10_21, data_operandA[11], data_operandB[10]);
	and stg_0_10_22(w_stg_0_10_22, data_operandA[12], data_operandB[10]);
	and stg_0_10_23(w_stg_0_10_23, data_operandA[13], data_operandB[10]);
	and stg_0_10_24(w_stg_0_10_24, data_operandA[14], data_operandB[10]);
	and stg_0_10_25(w_stg_0_10_25, data_operandA[15], data_operandB[10]);
	and stg_0_10_26(w_stg_0_10_26, data_operandA[16], data_operandB[10]);
	and stg_0_10_27(w_stg_0_10_27, data_operandA[17], data_operandB[10]);
	and stg_0_10_28(w_stg_0_10_28, data_operandA[18], data_operandB[10]);
	and stg_0_10_29(w_stg_0_10_29, data_operandA[19], data_operandB[10]);
	and stg_0_10_30(w_stg_0_10_30, data_operandA[20], data_operandB[10]);
	and stg_0_10_31(w_stg_0_10_31, data_operandA[21], data_operandB[10]);
	and stg_0_10_32(w_stg_0_10_32, data_operandA[22], data_operandB[10]);
	and stg_0_10_33(w_stg_0_10_33, data_operandA[23], data_operandB[10]);
	and stg_0_10_34(w_stg_0_10_34, data_operandA[24], data_operandB[10]);
	and stg_0_10_35(w_stg_0_10_35, data_operandA[25], data_operandB[10]);
	and stg_0_10_36(w_stg_0_10_36, data_operandA[26], data_operandB[10]);
	and stg_0_10_37(w_stg_0_10_37, data_operandA[27], data_operandB[10]);
	and stg_0_10_38(w_stg_0_10_38, data_operandA[28], data_operandB[10]);
	and stg_0_10_39(w_stg_0_10_39, data_operandA[29], data_operandB[10]);
	and stg_0_10_40(w_stg_0_10_40, data_operandA[30], data_operandB[10]);
	and stg_0_10_41(w_stg_0_10_41, data_operandA[31], data_operandB[10]);
	and stg_0_11_11(w_stg_0_11_11, data_operandA[0], data_operandB[11]);
	and stg_0_11_12(w_stg_0_11_12, data_operandA[1], data_operandB[11]);
	and stg_0_11_13(w_stg_0_11_13, data_operandA[2], data_operandB[11]);
	and stg_0_11_14(w_stg_0_11_14, data_operandA[3], data_operandB[11]);
	and stg_0_11_15(w_stg_0_11_15, data_operandA[4], data_operandB[11]);
	and stg_0_11_16(w_stg_0_11_16, data_operandA[5], data_operandB[11]);
	and stg_0_11_17(w_stg_0_11_17, data_operandA[6], data_operandB[11]);
	and stg_0_11_18(w_stg_0_11_18, data_operandA[7], data_operandB[11]);
	and stg_0_11_19(w_stg_0_11_19, data_operandA[8], data_operandB[11]);
	and stg_0_11_20(w_stg_0_11_20, data_operandA[9], data_operandB[11]);
	and stg_0_11_21(w_stg_0_11_21, data_operandA[10], data_operandB[11]);
	and stg_0_11_22(w_stg_0_11_22, data_operandA[11], data_operandB[11]);
	and stg_0_11_23(w_stg_0_11_23, data_operandA[12], data_operandB[11]);
	and stg_0_11_24(w_stg_0_11_24, data_operandA[13], data_operandB[11]);
	and stg_0_11_25(w_stg_0_11_25, data_operandA[14], data_operandB[11]);
	and stg_0_11_26(w_stg_0_11_26, data_operandA[15], data_operandB[11]);
	and stg_0_11_27(w_stg_0_11_27, data_operandA[16], data_operandB[11]);
	and stg_0_11_28(w_stg_0_11_28, data_operandA[17], data_operandB[11]);
	and stg_0_11_29(w_stg_0_11_29, data_operandA[18], data_operandB[11]);
	and stg_0_11_30(w_stg_0_11_30, data_operandA[19], data_operandB[11]);
	and stg_0_11_31(w_stg_0_11_31, data_operandA[20], data_operandB[11]);
	and stg_0_11_32(w_stg_0_11_32, data_operandA[21], data_operandB[11]);
	and stg_0_11_33(w_stg_0_11_33, data_operandA[22], data_operandB[11]);
	and stg_0_11_34(w_stg_0_11_34, data_operandA[23], data_operandB[11]);
	and stg_0_11_35(w_stg_0_11_35, data_operandA[24], data_operandB[11]);
	and stg_0_11_36(w_stg_0_11_36, data_operandA[25], data_operandB[11]);
	and stg_0_11_37(w_stg_0_11_37, data_operandA[26], data_operandB[11]);
	and stg_0_11_38(w_stg_0_11_38, data_operandA[27], data_operandB[11]);
	and stg_0_11_39(w_stg_0_11_39, data_operandA[28], data_operandB[11]);
	and stg_0_11_40(w_stg_0_11_40, data_operandA[29], data_operandB[11]);
	and stg_0_11_41(w_stg_0_11_41, data_operandA[30], data_operandB[11]);
	and stg_0_11_42(w_stg_0_11_42, data_operandA[31], data_operandB[11]);
	and stg_0_12_12(w_stg_0_12_12, data_operandA[0], data_operandB[12]);
	and stg_0_12_13(w_stg_0_12_13, data_operandA[1], data_operandB[12]);
	and stg_0_12_14(w_stg_0_12_14, data_operandA[2], data_operandB[12]);
	and stg_0_12_15(w_stg_0_12_15, data_operandA[3], data_operandB[12]);
	and stg_0_12_16(w_stg_0_12_16, data_operandA[4], data_operandB[12]);
	and stg_0_12_17(w_stg_0_12_17, data_operandA[5], data_operandB[12]);
	and stg_0_12_18(w_stg_0_12_18, data_operandA[6], data_operandB[12]);
	and stg_0_12_19(w_stg_0_12_19, data_operandA[7], data_operandB[12]);
	and stg_0_12_20(w_stg_0_12_20, data_operandA[8], data_operandB[12]);
	and stg_0_12_21(w_stg_0_12_21, data_operandA[9], data_operandB[12]);
	and stg_0_12_22(w_stg_0_12_22, data_operandA[10], data_operandB[12]);
	and stg_0_12_23(w_stg_0_12_23, data_operandA[11], data_operandB[12]);
	and stg_0_12_24(w_stg_0_12_24, data_operandA[12], data_operandB[12]);
	and stg_0_12_25(w_stg_0_12_25, data_operandA[13], data_operandB[12]);
	and stg_0_12_26(w_stg_0_12_26, data_operandA[14], data_operandB[12]);
	and stg_0_12_27(w_stg_0_12_27, data_operandA[15], data_operandB[12]);
	and stg_0_12_28(w_stg_0_12_28, data_operandA[16], data_operandB[12]);
	and stg_0_12_29(w_stg_0_12_29, data_operandA[17], data_operandB[12]);
	and stg_0_12_30(w_stg_0_12_30, data_operandA[18], data_operandB[12]);
	and stg_0_12_31(w_stg_0_12_31, data_operandA[19], data_operandB[12]);
	and stg_0_12_32(w_stg_0_12_32, data_operandA[20], data_operandB[12]);
	and stg_0_12_33(w_stg_0_12_33, data_operandA[21], data_operandB[12]);
	and stg_0_12_34(w_stg_0_12_34, data_operandA[22], data_operandB[12]);
	and stg_0_12_35(w_stg_0_12_35, data_operandA[23], data_operandB[12]);
	and stg_0_12_36(w_stg_0_12_36, data_operandA[24], data_operandB[12]);
	and stg_0_12_37(w_stg_0_12_37, data_operandA[25], data_operandB[12]);
	and stg_0_12_38(w_stg_0_12_38, data_operandA[26], data_operandB[12]);
	and stg_0_12_39(w_stg_0_12_39, data_operandA[27], data_operandB[12]);
	and stg_0_12_40(w_stg_0_12_40, data_operandA[28], data_operandB[12]);
	and stg_0_12_41(w_stg_0_12_41, data_operandA[29], data_operandB[12]);
	and stg_0_12_42(w_stg_0_12_42, data_operandA[30], data_operandB[12]);
	and stg_0_12_43(w_stg_0_12_43, data_operandA[31], data_operandB[12]);
	and stg_0_13_13(w_stg_0_13_13, data_operandA[0], data_operandB[13]);
	and stg_0_13_14(w_stg_0_13_14, data_operandA[1], data_operandB[13]);
	and stg_0_13_15(w_stg_0_13_15, data_operandA[2], data_operandB[13]);
	and stg_0_13_16(w_stg_0_13_16, data_operandA[3], data_operandB[13]);
	and stg_0_13_17(w_stg_0_13_17, data_operandA[4], data_operandB[13]);
	and stg_0_13_18(w_stg_0_13_18, data_operandA[5], data_operandB[13]);
	and stg_0_13_19(w_stg_0_13_19, data_operandA[6], data_operandB[13]);
	and stg_0_13_20(w_stg_0_13_20, data_operandA[7], data_operandB[13]);
	and stg_0_13_21(w_stg_0_13_21, data_operandA[8], data_operandB[13]);
	and stg_0_13_22(w_stg_0_13_22, data_operandA[9], data_operandB[13]);
	and stg_0_13_23(w_stg_0_13_23, data_operandA[10], data_operandB[13]);
	and stg_0_13_24(w_stg_0_13_24, data_operandA[11], data_operandB[13]);
	and stg_0_13_25(w_stg_0_13_25, data_operandA[12], data_operandB[13]);
	and stg_0_13_26(w_stg_0_13_26, data_operandA[13], data_operandB[13]);
	and stg_0_13_27(w_stg_0_13_27, data_operandA[14], data_operandB[13]);
	and stg_0_13_28(w_stg_0_13_28, data_operandA[15], data_operandB[13]);
	and stg_0_13_29(w_stg_0_13_29, data_operandA[16], data_operandB[13]);
	and stg_0_13_30(w_stg_0_13_30, data_operandA[17], data_operandB[13]);
	and stg_0_13_31(w_stg_0_13_31, data_operandA[18], data_operandB[13]);
	and stg_0_13_32(w_stg_0_13_32, data_operandA[19], data_operandB[13]);
	and stg_0_13_33(w_stg_0_13_33, data_operandA[20], data_operandB[13]);
	and stg_0_13_34(w_stg_0_13_34, data_operandA[21], data_operandB[13]);
	and stg_0_13_35(w_stg_0_13_35, data_operandA[22], data_operandB[13]);
	and stg_0_13_36(w_stg_0_13_36, data_operandA[23], data_operandB[13]);
	and stg_0_13_37(w_stg_0_13_37, data_operandA[24], data_operandB[13]);
	and stg_0_13_38(w_stg_0_13_38, data_operandA[25], data_operandB[13]);
	and stg_0_13_39(w_stg_0_13_39, data_operandA[26], data_operandB[13]);
	and stg_0_13_40(w_stg_0_13_40, data_operandA[27], data_operandB[13]);
	and stg_0_13_41(w_stg_0_13_41, data_operandA[28], data_operandB[13]);
	and stg_0_13_42(w_stg_0_13_42, data_operandA[29], data_operandB[13]);
	and stg_0_13_43(w_stg_0_13_43, data_operandA[30], data_operandB[13]);
	and stg_0_13_44(w_stg_0_13_44, data_operandA[31], data_operandB[13]);
	and stg_0_14_14(w_stg_0_14_14, data_operandA[0], data_operandB[14]);
	and stg_0_14_15(w_stg_0_14_15, data_operandA[1], data_operandB[14]);
	and stg_0_14_16(w_stg_0_14_16, data_operandA[2], data_operandB[14]);
	and stg_0_14_17(w_stg_0_14_17, data_operandA[3], data_operandB[14]);
	and stg_0_14_18(w_stg_0_14_18, data_operandA[4], data_operandB[14]);
	and stg_0_14_19(w_stg_0_14_19, data_operandA[5], data_operandB[14]);
	and stg_0_14_20(w_stg_0_14_20, data_operandA[6], data_operandB[14]);
	and stg_0_14_21(w_stg_0_14_21, data_operandA[7], data_operandB[14]);
	and stg_0_14_22(w_stg_0_14_22, data_operandA[8], data_operandB[14]);
	and stg_0_14_23(w_stg_0_14_23, data_operandA[9], data_operandB[14]);
	and stg_0_14_24(w_stg_0_14_24, data_operandA[10], data_operandB[14]);
	and stg_0_14_25(w_stg_0_14_25, data_operandA[11], data_operandB[14]);
	and stg_0_14_26(w_stg_0_14_26, data_operandA[12], data_operandB[14]);
	and stg_0_14_27(w_stg_0_14_27, data_operandA[13], data_operandB[14]);
	and stg_0_14_28(w_stg_0_14_28, data_operandA[14], data_operandB[14]);
	and stg_0_14_29(w_stg_0_14_29, data_operandA[15], data_operandB[14]);
	and stg_0_14_30(w_stg_0_14_30, data_operandA[16], data_operandB[14]);
	and stg_0_14_31(w_stg_0_14_31, data_operandA[17], data_operandB[14]);
	and stg_0_14_32(w_stg_0_14_32, data_operandA[18], data_operandB[14]);
	and stg_0_14_33(w_stg_0_14_33, data_operandA[19], data_operandB[14]);
	and stg_0_14_34(w_stg_0_14_34, data_operandA[20], data_operandB[14]);
	and stg_0_14_35(w_stg_0_14_35, data_operandA[21], data_operandB[14]);
	and stg_0_14_36(w_stg_0_14_36, data_operandA[22], data_operandB[14]);
	and stg_0_14_37(w_stg_0_14_37, data_operandA[23], data_operandB[14]);
	and stg_0_14_38(w_stg_0_14_38, data_operandA[24], data_operandB[14]);
	and stg_0_14_39(w_stg_0_14_39, data_operandA[25], data_operandB[14]);
	and stg_0_14_40(w_stg_0_14_40, data_operandA[26], data_operandB[14]);
	and stg_0_14_41(w_stg_0_14_41, data_operandA[27], data_operandB[14]);
	and stg_0_14_42(w_stg_0_14_42, data_operandA[28], data_operandB[14]);
	and stg_0_14_43(w_stg_0_14_43, data_operandA[29], data_operandB[14]);
	and stg_0_14_44(w_stg_0_14_44, data_operandA[30], data_operandB[14]);
	and stg_0_14_45(w_stg_0_14_45, data_operandA[31], data_operandB[14]);
	and stg_0_15_15(w_stg_0_15_15, data_operandA[0], data_operandB[15]);
	and stg_0_15_16(w_stg_0_15_16, data_operandA[1], data_operandB[15]);
	and stg_0_15_17(w_stg_0_15_17, data_operandA[2], data_operandB[15]);
	and stg_0_15_18(w_stg_0_15_18, data_operandA[3], data_operandB[15]);
	and stg_0_15_19(w_stg_0_15_19, data_operandA[4], data_operandB[15]);
	and stg_0_15_20(w_stg_0_15_20, data_operandA[5], data_operandB[15]);
	and stg_0_15_21(w_stg_0_15_21, data_operandA[6], data_operandB[15]);
	and stg_0_15_22(w_stg_0_15_22, data_operandA[7], data_operandB[15]);
	and stg_0_15_23(w_stg_0_15_23, data_operandA[8], data_operandB[15]);
	and stg_0_15_24(w_stg_0_15_24, data_operandA[9], data_operandB[15]);
	and stg_0_15_25(w_stg_0_15_25, data_operandA[10], data_operandB[15]);
	and stg_0_15_26(w_stg_0_15_26, data_operandA[11], data_operandB[15]);
	and stg_0_15_27(w_stg_0_15_27, data_operandA[12], data_operandB[15]);
	and stg_0_15_28(w_stg_0_15_28, data_operandA[13], data_operandB[15]);
	and stg_0_15_29(w_stg_0_15_29, data_operandA[14], data_operandB[15]);
	and stg_0_15_30(w_stg_0_15_30, data_operandA[15], data_operandB[15]);
	and stg_0_15_31(w_stg_0_15_31, data_operandA[16], data_operandB[15]);
	and stg_0_15_32(w_stg_0_15_32, data_operandA[17], data_operandB[15]);
	and stg_0_15_33(w_stg_0_15_33, data_operandA[18], data_operandB[15]);
	and stg_0_15_34(w_stg_0_15_34, data_operandA[19], data_operandB[15]);
	and stg_0_15_35(w_stg_0_15_35, data_operandA[20], data_operandB[15]);
	and stg_0_15_36(w_stg_0_15_36, data_operandA[21], data_operandB[15]);
	and stg_0_15_37(w_stg_0_15_37, data_operandA[22], data_operandB[15]);
	and stg_0_15_38(w_stg_0_15_38, data_operandA[23], data_operandB[15]);
	and stg_0_15_39(w_stg_0_15_39, data_operandA[24], data_operandB[15]);
	and stg_0_15_40(w_stg_0_15_40, data_operandA[25], data_operandB[15]);
	and stg_0_15_41(w_stg_0_15_41, data_operandA[26], data_operandB[15]);
	and stg_0_15_42(w_stg_0_15_42, data_operandA[27], data_operandB[15]);
	and stg_0_15_43(w_stg_0_15_43, data_operandA[28], data_operandB[15]);
	and stg_0_15_44(w_stg_0_15_44, data_operandA[29], data_operandB[15]);
	and stg_0_15_45(w_stg_0_15_45, data_operandA[30], data_operandB[15]);
	and stg_0_15_46(w_stg_0_15_46, data_operandA[31], data_operandB[15]);
	and stg_0_16_16(w_stg_0_16_16, data_operandA[0], data_operandB[16]);
	and stg_0_16_17(w_stg_0_16_17, data_operandA[1], data_operandB[16]);
	and stg_0_16_18(w_stg_0_16_18, data_operandA[2], data_operandB[16]);
	and stg_0_16_19(w_stg_0_16_19, data_operandA[3], data_operandB[16]);
	and stg_0_16_20(w_stg_0_16_20, data_operandA[4], data_operandB[16]);
	and stg_0_16_21(w_stg_0_16_21, data_operandA[5], data_operandB[16]);
	and stg_0_16_22(w_stg_0_16_22, data_operandA[6], data_operandB[16]);
	and stg_0_16_23(w_stg_0_16_23, data_operandA[7], data_operandB[16]);
	and stg_0_16_24(w_stg_0_16_24, data_operandA[8], data_operandB[16]);
	and stg_0_16_25(w_stg_0_16_25, data_operandA[9], data_operandB[16]);
	and stg_0_16_26(w_stg_0_16_26, data_operandA[10], data_operandB[16]);
	and stg_0_16_27(w_stg_0_16_27, data_operandA[11], data_operandB[16]);
	and stg_0_16_28(w_stg_0_16_28, data_operandA[12], data_operandB[16]);
	and stg_0_16_29(w_stg_0_16_29, data_operandA[13], data_operandB[16]);
	and stg_0_16_30(w_stg_0_16_30, data_operandA[14], data_operandB[16]);
	and stg_0_16_31(w_stg_0_16_31, data_operandA[15], data_operandB[16]);
	and stg_0_16_32(w_stg_0_16_32, data_operandA[16], data_operandB[16]);
	and stg_0_16_33(w_stg_0_16_33, data_operandA[17], data_operandB[16]);
	and stg_0_16_34(w_stg_0_16_34, data_operandA[18], data_operandB[16]);
	and stg_0_16_35(w_stg_0_16_35, data_operandA[19], data_operandB[16]);
	and stg_0_16_36(w_stg_0_16_36, data_operandA[20], data_operandB[16]);
	and stg_0_16_37(w_stg_0_16_37, data_operandA[21], data_operandB[16]);
	and stg_0_16_38(w_stg_0_16_38, data_operandA[22], data_operandB[16]);
	and stg_0_16_39(w_stg_0_16_39, data_operandA[23], data_operandB[16]);
	and stg_0_16_40(w_stg_0_16_40, data_operandA[24], data_operandB[16]);
	and stg_0_16_41(w_stg_0_16_41, data_operandA[25], data_operandB[16]);
	and stg_0_16_42(w_stg_0_16_42, data_operandA[26], data_operandB[16]);
	and stg_0_16_43(w_stg_0_16_43, data_operandA[27], data_operandB[16]);
	and stg_0_16_44(w_stg_0_16_44, data_operandA[28], data_operandB[16]);
	and stg_0_16_45(w_stg_0_16_45, data_operandA[29], data_operandB[16]);
	and stg_0_16_46(w_stg_0_16_46, data_operandA[30], data_operandB[16]);
	and stg_0_16_47(w_stg_0_16_47, data_operandA[31], data_operandB[16]);
	and stg_0_17_17(w_stg_0_17_17, data_operandA[0], data_operandB[17]);
	and stg_0_17_18(w_stg_0_17_18, data_operandA[1], data_operandB[17]);
	and stg_0_17_19(w_stg_0_17_19, data_operandA[2], data_operandB[17]);
	and stg_0_17_20(w_stg_0_17_20, data_operandA[3], data_operandB[17]);
	and stg_0_17_21(w_stg_0_17_21, data_operandA[4], data_operandB[17]);
	and stg_0_17_22(w_stg_0_17_22, data_operandA[5], data_operandB[17]);
	and stg_0_17_23(w_stg_0_17_23, data_operandA[6], data_operandB[17]);
	and stg_0_17_24(w_stg_0_17_24, data_operandA[7], data_operandB[17]);
	and stg_0_17_25(w_stg_0_17_25, data_operandA[8], data_operandB[17]);
	and stg_0_17_26(w_stg_0_17_26, data_operandA[9], data_operandB[17]);
	and stg_0_17_27(w_stg_0_17_27, data_operandA[10], data_operandB[17]);
	and stg_0_17_28(w_stg_0_17_28, data_operandA[11], data_operandB[17]);
	and stg_0_17_29(w_stg_0_17_29, data_operandA[12], data_operandB[17]);
	and stg_0_17_30(w_stg_0_17_30, data_operandA[13], data_operandB[17]);
	and stg_0_17_31(w_stg_0_17_31, data_operandA[14], data_operandB[17]);
	and stg_0_17_32(w_stg_0_17_32, data_operandA[15], data_operandB[17]);
	and stg_0_17_33(w_stg_0_17_33, data_operandA[16], data_operandB[17]);
	and stg_0_17_34(w_stg_0_17_34, data_operandA[17], data_operandB[17]);
	and stg_0_17_35(w_stg_0_17_35, data_operandA[18], data_operandB[17]);
	and stg_0_17_36(w_stg_0_17_36, data_operandA[19], data_operandB[17]);
	and stg_0_17_37(w_stg_0_17_37, data_operandA[20], data_operandB[17]);
	and stg_0_17_38(w_stg_0_17_38, data_operandA[21], data_operandB[17]);
	and stg_0_17_39(w_stg_0_17_39, data_operandA[22], data_operandB[17]);
	and stg_0_17_40(w_stg_0_17_40, data_operandA[23], data_operandB[17]);
	and stg_0_17_41(w_stg_0_17_41, data_operandA[24], data_operandB[17]);
	and stg_0_17_42(w_stg_0_17_42, data_operandA[25], data_operandB[17]);
	and stg_0_17_43(w_stg_0_17_43, data_operandA[26], data_operandB[17]);
	and stg_0_17_44(w_stg_0_17_44, data_operandA[27], data_operandB[17]);
	and stg_0_17_45(w_stg_0_17_45, data_operandA[28], data_operandB[17]);
	and stg_0_17_46(w_stg_0_17_46, data_operandA[29], data_operandB[17]);
	and stg_0_17_47(w_stg_0_17_47, data_operandA[30], data_operandB[17]);
	and stg_0_17_48(w_stg_0_17_48, data_operandA[31], data_operandB[17]);
	and stg_0_18_18(w_stg_0_18_18, data_operandA[0], data_operandB[18]);
	and stg_0_18_19(w_stg_0_18_19, data_operandA[1], data_operandB[18]);
	and stg_0_18_20(w_stg_0_18_20, data_operandA[2], data_operandB[18]);
	and stg_0_18_21(w_stg_0_18_21, data_operandA[3], data_operandB[18]);
	and stg_0_18_22(w_stg_0_18_22, data_operandA[4], data_operandB[18]);
	and stg_0_18_23(w_stg_0_18_23, data_operandA[5], data_operandB[18]);
	and stg_0_18_24(w_stg_0_18_24, data_operandA[6], data_operandB[18]);
	and stg_0_18_25(w_stg_0_18_25, data_operandA[7], data_operandB[18]);
	and stg_0_18_26(w_stg_0_18_26, data_operandA[8], data_operandB[18]);
	and stg_0_18_27(w_stg_0_18_27, data_operandA[9], data_operandB[18]);
	and stg_0_18_28(w_stg_0_18_28, data_operandA[10], data_operandB[18]);
	and stg_0_18_29(w_stg_0_18_29, data_operandA[11], data_operandB[18]);
	and stg_0_18_30(w_stg_0_18_30, data_operandA[12], data_operandB[18]);
	and stg_0_18_31(w_stg_0_18_31, data_operandA[13], data_operandB[18]);
	and stg_0_18_32(w_stg_0_18_32, data_operandA[14], data_operandB[18]);
	and stg_0_18_33(w_stg_0_18_33, data_operandA[15], data_operandB[18]);
	and stg_0_18_34(w_stg_0_18_34, data_operandA[16], data_operandB[18]);
	and stg_0_18_35(w_stg_0_18_35, data_operandA[17], data_operandB[18]);
	and stg_0_18_36(w_stg_0_18_36, data_operandA[18], data_operandB[18]);
	and stg_0_18_37(w_stg_0_18_37, data_operandA[19], data_operandB[18]);
	and stg_0_18_38(w_stg_0_18_38, data_operandA[20], data_operandB[18]);
	and stg_0_18_39(w_stg_0_18_39, data_operandA[21], data_operandB[18]);
	and stg_0_18_40(w_stg_0_18_40, data_operandA[22], data_operandB[18]);
	and stg_0_18_41(w_stg_0_18_41, data_operandA[23], data_operandB[18]);
	and stg_0_18_42(w_stg_0_18_42, data_operandA[24], data_operandB[18]);
	and stg_0_18_43(w_stg_0_18_43, data_operandA[25], data_operandB[18]);
	and stg_0_18_44(w_stg_0_18_44, data_operandA[26], data_operandB[18]);
	and stg_0_18_45(w_stg_0_18_45, data_operandA[27], data_operandB[18]);
	and stg_0_18_46(w_stg_0_18_46, data_operandA[28], data_operandB[18]);
	and stg_0_18_47(w_stg_0_18_47, data_operandA[29], data_operandB[18]);
	and stg_0_18_48(w_stg_0_18_48, data_operandA[30], data_operandB[18]);
	and stg_0_18_49(w_stg_0_18_49, data_operandA[31], data_operandB[18]);
	and stg_0_19_19(w_stg_0_19_19, data_operandA[0], data_operandB[19]);
	and stg_0_19_20(w_stg_0_19_20, data_operandA[1], data_operandB[19]);
	and stg_0_19_21(w_stg_0_19_21, data_operandA[2], data_operandB[19]);
	and stg_0_19_22(w_stg_0_19_22, data_operandA[3], data_operandB[19]);
	and stg_0_19_23(w_stg_0_19_23, data_operandA[4], data_operandB[19]);
	and stg_0_19_24(w_stg_0_19_24, data_operandA[5], data_operandB[19]);
	and stg_0_19_25(w_stg_0_19_25, data_operandA[6], data_operandB[19]);
	and stg_0_19_26(w_stg_0_19_26, data_operandA[7], data_operandB[19]);
	and stg_0_19_27(w_stg_0_19_27, data_operandA[8], data_operandB[19]);
	and stg_0_19_28(w_stg_0_19_28, data_operandA[9], data_operandB[19]);
	and stg_0_19_29(w_stg_0_19_29, data_operandA[10], data_operandB[19]);
	and stg_0_19_30(w_stg_0_19_30, data_operandA[11], data_operandB[19]);
	and stg_0_19_31(w_stg_0_19_31, data_operandA[12], data_operandB[19]);
	and stg_0_19_32(w_stg_0_19_32, data_operandA[13], data_operandB[19]);
	and stg_0_19_33(w_stg_0_19_33, data_operandA[14], data_operandB[19]);
	and stg_0_19_34(w_stg_0_19_34, data_operandA[15], data_operandB[19]);
	and stg_0_19_35(w_stg_0_19_35, data_operandA[16], data_operandB[19]);
	and stg_0_19_36(w_stg_0_19_36, data_operandA[17], data_operandB[19]);
	and stg_0_19_37(w_stg_0_19_37, data_operandA[18], data_operandB[19]);
	and stg_0_19_38(w_stg_0_19_38, data_operandA[19], data_operandB[19]);
	and stg_0_19_39(w_stg_0_19_39, data_operandA[20], data_operandB[19]);
	and stg_0_19_40(w_stg_0_19_40, data_operandA[21], data_operandB[19]);
	and stg_0_19_41(w_stg_0_19_41, data_operandA[22], data_operandB[19]);
	and stg_0_19_42(w_stg_0_19_42, data_operandA[23], data_operandB[19]);
	and stg_0_19_43(w_stg_0_19_43, data_operandA[24], data_operandB[19]);
	and stg_0_19_44(w_stg_0_19_44, data_operandA[25], data_operandB[19]);
	and stg_0_19_45(w_stg_0_19_45, data_operandA[26], data_operandB[19]);
	and stg_0_19_46(w_stg_0_19_46, data_operandA[27], data_operandB[19]);
	and stg_0_19_47(w_stg_0_19_47, data_operandA[28], data_operandB[19]);
	and stg_0_19_48(w_stg_0_19_48, data_operandA[29], data_operandB[19]);
	and stg_0_19_49(w_stg_0_19_49, data_operandA[30], data_operandB[19]);
	and stg_0_19_50(w_stg_0_19_50, data_operandA[31], data_operandB[19]);
	and stg_0_20_20(w_stg_0_20_20, data_operandA[0], data_operandB[20]);
	and stg_0_20_21(w_stg_0_20_21, data_operandA[1], data_operandB[20]);
	and stg_0_20_22(w_stg_0_20_22, data_operandA[2], data_operandB[20]);
	and stg_0_20_23(w_stg_0_20_23, data_operandA[3], data_operandB[20]);
	and stg_0_20_24(w_stg_0_20_24, data_operandA[4], data_operandB[20]);
	and stg_0_20_25(w_stg_0_20_25, data_operandA[5], data_operandB[20]);
	and stg_0_20_26(w_stg_0_20_26, data_operandA[6], data_operandB[20]);
	and stg_0_20_27(w_stg_0_20_27, data_operandA[7], data_operandB[20]);
	and stg_0_20_28(w_stg_0_20_28, data_operandA[8], data_operandB[20]);
	and stg_0_20_29(w_stg_0_20_29, data_operandA[9], data_operandB[20]);
	and stg_0_20_30(w_stg_0_20_30, data_operandA[10], data_operandB[20]);
	and stg_0_20_31(w_stg_0_20_31, data_operandA[11], data_operandB[20]);
	and stg_0_20_32(w_stg_0_20_32, data_operandA[12], data_operandB[20]);
	and stg_0_20_33(w_stg_0_20_33, data_operandA[13], data_operandB[20]);
	and stg_0_20_34(w_stg_0_20_34, data_operandA[14], data_operandB[20]);
	and stg_0_20_35(w_stg_0_20_35, data_operandA[15], data_operandB[20]);
	and stg_0_20_36(w_stg_0_20_36, data_operandA[16], data_operandB[20]);
	and stg_0_20_37(w_stg_0_20_37, data_operandA[17], data_operandB[20]);
	and stg_0_20_38(w_stg_0_20_38, data_operandA[18], data_operandB[20]);
	and stg_0_20_39(w_stg_0_20_39, data_operandA[19], data_operandB[20]);
	and stg_0_20_40(w_stg_0_20_40, data_operandA[20], data_operandB[20]);
	and stg_0_20_41(w_stg_0_20_41, data_operandA[21], data_operandB[20]);
	and stg_0_20_42(w_stg_0_20_42, data_operandA[22], data_operandB[20]);
	and stg_0_20_43(w_stg_0_20_43, data_operandA[23], data_operandB[20]);
	and stg_0_20_44(w_stg_0_20_44, data_operandA[24], data_operandB[20]);
	and stg_0_20_45(w_stg_0_20_45, data_operandA[25], data_operandB[20]);
	and stg_0_20_46(w_stg_0_20_46, data_operandA[26], data_operandB[20]);
	and stg_0_20_47(w_stg_0_20_47, data_operandA[27], data_operandB[20]);
	and stg_0_20_48(w_stg_0_20_48, data_operandA[28], data_operandB[20]);
	and stg_0_20_49(w_stg_0_20_49, data_operandA[29], data_operandB[20]);
	and stg_0_20_50(w_stg_0_20_50, data_operandA[30], data_operandB[20]);
	and stg_0_20_51(w_stg_0_20_51, data_operandA[31], data_operandB[20]);
	and stg_0_21_21(w_stg_0_21_21, data_operandA[0], data_operandB[21]);
	and stg_0_21_22(w_stg_0_21_22, data_operandA[1], data_operandB[21]);
	and stg_0_21_23(w_stg_0_21_23, data_operandA[2], data_operandB[21]);
	and stg_0_21_24(w_stg_0_21_24, data_operandA[3], data_operandB[21]);
	and stg_0_21_25(w_stg_0_21_25, data_operandA[4], data_operandB[21]);
	and stg_0_21_26(w_stg_0_21_26, data_operandA[5], data_operandB[21]);
	and stg_0_21_27(w_stg_0_21_27, data_operandA[6], data_operandB[21]);
	and stg_0_21_28(w_stg_0_21_28, data_operandA[7], data_operandB[21]);
	and stg_0_21_29(w_stg_0_21_29, data_operandA[8], data_operandB[21]);
	and stg_0_21_30(w_stg_0_21_30, data_operandA[9], data_operandB[21]);
	and stg_0_21_31(w_stg_0_21_31, data_operandA[10], data_operandB[21]);
	and stg_0_21_32(w_stg_0_21_32, data_operandA[11], data_operandB[21]);
	and stg_0_21_33(w_stg_0_21_33, data_operandA[12], data_operandB[21]);
	and stg_0_21_34(w_stg_0_21_34, data_operandA[13], data_operandB[21]);
	and stg_0_21_35(w_stg_0_21_35, data_operandA[14], data_operandB[21]);
	and stg_0_21_36(w_stg_0_21_36, data_operandA[15], data_operandB[21]);
	and stg_0_21_37(w_stg_0_21_37, data_operandA[16], data_operandB[21]);
	and stg_0_21_38(w_stg_0_21_38, data_operandA[17], data_operandB[21]);
	and stg_0_21_39(w_stg_0_21_39, data_operandA[18], data_operandB[21]);
	and stg_0_21_40(w_stg_0_21_40, data_operandA[19], data_operandB[21]);
	and stg_0_21_41(w_stg_0_21_41, data_operandA[20], data_operandB[21]);
	and stg_0_21_42(w_stg_0_21_42, data_operandA[21], data_operandB[21]);
	and stg_0_21_43(w_stg_0_21_43, data_operandA[22], data_operandB[21]);
	and stg_0_21_44(w_stg_0_21_44, data_operandA[23], data_operandB[21]);
	and stg_0_21_45(w_stg_0_21_45, data_operandA[24], data_operandB[21]);
	and stg_0_21_46(w_stg_0_21_46, data_operandA[25], data_operandB[21]);
	and stg_0_21_47(w_stg_0_21_47, data_operandA[26], data_operandB[21]);
	and stg_0_21_48(w_stg_0_21_48, data_operandA[27], data_operandB[21]);
	and stg_0_21_49(w_stg_0_21_49, data_operandA[28], data_operandB[21]);
	and stg_0_21_50(w_stg_0_21_50, data_operandA[29], data_operandB[21]);
	and stg_0_21_51(w_stg_0_21_51, data_operandA[30], data_operandB[21]);
	and stg_0_21_52(w_stg_0_21_52, data_operandA[31], data_operandB[21]);
	and stg_0_22_22(w_stg_0_22_22, data_operandA[0], data_operandB[22]);
	and stg_0_22_23(w_stg_0_22_23, data_operandA[1], data_operandB[22]);
	and stg_0_22_24(w_stg_0_22_24, data_operandA[2], data_operandB[22]);
	and stg_0_22_25(w_stg_0_22_25, data_operandA[3], data_operandB[22]);
	and stg_0_22_26(w_stg_0_22_26, data_operandA[4], data_operandB[22]);
	and stg_0_22_27(w_stg_0_22_27, data_operandA[5], data_operandB[22]);
	and stg_0_22_28(w_stg_0_22_28, data_operandA[6], data_operandB[22]);
	and stg_0_22_29(w_stg_0_22_29, data_operandA[7], data_operandB[22]);
	and stg_0_22_30(w_stg_0_22_30, data_operandA[8], data_operandB[22]);
	and stg_0_22_31(w_stg_0_22_31, data_operandA[9], data_operandB[22]);
	and stg_0_22_32(w_stg_0_22_32, data_operandA[10], data_operandB[22]);
	and stg_0_22_33(w_stg_0_22_33, data_operandA[11], data_operandB[22]);
	and stg_0_22_34(w_stg_0_22_34, data_operandA[12], data_operandB[22]);
	and stg_0_22_35(w_stg_0_22_35, data_operandA[13], data_operandB[22]);
	and stg_0_22_36(w_stg_0_22_36, data_operandA[14], data_operandB[22]);
	and stg_0_22_37(w_stg_0_22_37, data_operandA[15], data_operandB[22]);
	and stg_0_22_38(w_stg_0_22_38, data_operandA[16], data_operandB[22]);
	and stg_0_22_39(w_stg_0_22_39, data_operandA[17], data_operandB[22]);
	and stg_0_22_40(w_stg_0_22_40, data_operandA[18], data_operandB[22]);
	and stg_0_22_41(w_stg_0_22_41, data_operandA[19], data_operandB[22]);
	and stg_0_22_42(w_stg_0_22_42, data_operandA[20], data_operandB[22]);
	and stg_0_22_43(w_stg_0_22_43, data_operandA[21], data_operandB[22]);
	and stg_0_22_44(w_stg_0_22_44, data_operandA[22], data_operandB[22]);
	and stg_0_22_45(w_stg_0_22_45, data_operandA[23], data_operandB[22]);
	and stg_0_22_46(w_stg_0_22_46, data_operandA[24], data_operandB[22]);
	and stg_0_22_47(w_stg_0_22_47, data_operandA[25], data_operandB[22]);
	and stg_0_22_48(w_stg_0_22_48, data_operandA[26], data_operandB[22]);
	and stg_0_22_49(w_stg_0_22_49, data_operandA[27], data_operandB[22]);
	and stg_0_22_50(w_stg_0_22_50, data_operandA[28], data_operandB[22]);
	and stg_0_22_51(w_stg_0_22_51, data_operandA[29], data_operandB[22]);
	and stg_0_22_52(w_stg_0_22_52, data_operandA[30], data_operandB[22]);
	and stg_0_22_53(w_stg_0_22_53, data_operandA[31], data_operandB[22]);
	and stg_0_23_23(w_stg_0_23_23, data_operandA[0], data_operandB[23]);
	and stg_0_23_24(w_stg_0_23_24, data_operandA[1], data_operandB[23]);
	and stg_0_23_25(w_stg_0_23_25, data_operandA[2], data_operandB[23]);
	and stg_0_23_26(w_stg_0_23_26, data_operandA[3], data_operandB[23]);
	and stg_0_23_27(w_stg_0_23_27, data_operandA[4], data_operandB[23]);
	and stg_0_23_28(w_stg_0_23_28, data_operandA[5], data_operandB[23]);
	and stg_0_23_29(w_stg_0_23_29, data_operandA[6], data_operandB[23]);
	and stg_0_23_30(w_stg_0_23_30, data_operandA[7], data_operandB[23]);
	and stg_0_23_31(w_stg_0_23_31, data_operandA[8], data_operandB[23]);
	and stg_0_23_32(w_stg_0_23_32, data_operandA[9], data_operandB[23]);
	and stg_0_23_33(w_stg_0_23_33, data_operandA[10], data_operandB[23]);
	and stg_0_23_34(w_stg_0_23_34, data_operandA[11], data_operandB[23]);
	and stg_0_23_35(w_stg_0_23_35, data_operandA[12], data_operandB[23]);
	and stg_0_23_36(w_stg_0_23_36, data_operandA[13], data_operandB[23]);
	and stg_0_23_37(w_stg_0_23_37, data_operandA[14], data_operandB[23]);
	and stg_0_23_38(w_stg_0_23_38, data_operandA[15], data_operandB[23]);
	and stg_0_23_39(w_stg_0_23_39, data_operandA[16], data_operandB[23]);
	and stg_0_23_40(w_stg_0_23_40, data_operandA[17], data_operandB[23]);
	and stg_0_23_41(w_stg_0_23_41, data_operandA[18], data_operandB[23]);
	and stg_0_23_42(w_stg_0_23_42, data_operandA[19], data_operandB[23]);
	and stg_0_23_43(w_stg_0_23_43, data_operandA[20], data_operandB[23]);
	and stg_0_23_44(w_stg_0_23_44, data_operandA[21], data_operandB[23]);
	and stg_0_23_45(w_stg_0_23_45, data_operandA[22], data_operandB[23]);
	and stg_0_23_46(w_stg_0_23_46, data_operandA[23], data_operandB[23]);
	and stg_0_23_47(w_stg_0_23_47, data_operandA[24], data_operandB[23]);
	and stg_0_23_48(w_stg_0_23_48, data_operandA[25], data_operandB[23]);
	and stg_0_23_49(w_stg_0_23_49, data_operandA[26], data_operandB[23]);
	and stg_0_23_50(w_stg_0_23_50, data_operandA[27], data_operandB[23]);
	and stg_0_23_51(w_stg_0_23_51, data_operandA[28], data_operandB[23]);
	and stg_0_23_52(w_stg_0_23_52, data_operandA[29], data_operandB[23]);
	and stg_0_23_53(w_stg_0_23_53, data_operandA[30], data_operandB[23]);
	and stg_0_23_54(w_stg_0_23_54, data_operandA[31], data_operandB[23]);
	and stg_0_24_24(w_stg_0_24_24, data_operandA[0], data_operandB[24]);
	and stg_0_24_25(w_stg_0_24_25, data_operandA[1], data_operandB[24]);
	and stg_0_24_26(w_stg_0_24_26, data_operandA[2], data_operandB[24]);
	and stg_0_24_27(w_stg_0_24_27, data_operandA[3], data_operandB[24]);
	and stg_0_24_28(w_stg_0_24_28, data_operandA[4], data_operandB[24]);
	and stg_0_24_29(w_stg_0_24_29, data_operandA[5], data_operandB[24]);
	and stg_0_24_30(w_stg_0_24_30, data_operandA[6], data_operandB[24]);
	and stg_0_24_31(w_stg_0_24_31, data_operandA[7], data_operandB[24]);
	and stg_0_24_32(w_stg_0_24_32, data_operandA[8], data_operandB[24]);
	and stg_0_24_33(w_stg_0_24_33, data_operandA[9], data_operandB[24]);
	and stg_0_24_34(w_stg_0_24_34, data_operandA[10], data_operandB[24]);
	and stg_0_24_35(w_stg_0_24_35, data_operandA[11], data_operandB[24]);
	and stg_0_24_36(w_stg_0_24_36, data_operandA[12], data_operandB[24]);
	and stg_0_24_37(w_stg_0_24_37, data_operandA[13], data_operandB[24]);
	and stg_0_24_38(w_stg_0_24_38, data_operandA[14], data_operandB[24]);
	and stg_0_24_39(w_stg_0_24_39, data_operandA[15], data_operandB[24]);
	and stg_0_24_40(w_stg_0_24_40, data_operandA[16], data_operandB[24]);
	and stg_0_24_41(w_stg_0_24_41, data_operandA[17], data_operandB[24]);
	and stg_0_24_42(w_stg_0_24_42, data_operandA[18], data_operandB[24]);
	and stg_0_24_43(w_stg_0_24_43, data_operandA[19], data_operandB[24]);
	and stg_0_24_44(w_stg_0_24_44, data_operandA[20], data_operandB[24]);
	and stg_0_24_45(w_stg_0_24_45, data_operandA[21], data_operandB[24]);
	and stg_0_24_46(w_stg_0_24_46, data_operandA[22], data_operandB[24]);
	and stg_0_24_47(w_stg_0_24_47, data_operandA[23], data_operandB[24]);
	and stg_0_24_48(w_stg_0_24_48, data_operandA[24], data_operandB[24]);
	and stg_0_24_49(w_stg_0_24_49, data_operandA[25], data_operandB[24]);
	and stg_0_24_50(w_stg_0_24_50, data_operandA[26], data_operandB[24]);
	and stg_0_24_51(w_stg_0_24_51, data_operandA[27], data_operandB[24]);
	and stg_0_24_52(w_stg_0_24_52, data_operandA[28], data_operandB[24]);
	and stg_0_24_53(w_stg_0_24_53, data_operandA[29], data_operandB[24]);
	and stg_0_24_54(w_stg_0_24_54, data_operandA[30], data_operandB[24]);
	and stg_0_24_55(w_stg_0_24_55, data_operandA[31], data_operandB[24]);
	and stg_0_25_25(w_stg_0_25_25, data_operandA[0], data_operandB[25]);
	and stg_0_25_26(w_stg_0_25_26, data_operandA[1], data_operandB[25]);
	and stg_0_25_27(w_stg_0_25_27, data_operandA[2], data_operandB[25]);
	and stg_0_25_28(w_stg_0_25_28, data_operandA[3], data_operandB[25]);
	and stg_0_25_29(w_stg_0_25_29, data_operandA[4], data_operandB[25]);
	and stg_0_25_30(w_stg_0_25_30, data_operandA[5], data_operandB[25]);
	and stg_0_25_31(w_stg_0_25_31, data_operandA[6], data_operandB[25]);
	and stg_0_25_32(w_stg_0_25_32, data_operandA[7], data_operandB[25]);
	and stg_0_25_33(w_stg_0_25_33, data_operandA[8], data_operandB[25]);
	and stg_0_25_34(w_stg_0_25_34, data_operandA[9], data_operandB[25]);
	and stg_0_25_35(w_stg_0_25_35, data_operandA[10], data_operandB[25]);
	and stg_0_25_36(w_stg_0_25_36, data_operandA[11], data_operandB[25]);
	and stg_0_25_37(w_stg_0_25_37, data_operandA[12], data_operandB[25]);
	and stg_0_25_38(w_stg_0_25_38, data_operandA[13], data_operandB[25]);
	and stg_0_25_39(w_stg_0_25_39, data_operandA[14], data_operandB[25]);
	and stg_0_25_40(w_stg_0_25_40, data_operandA[15], data_operandB[25]);
	and stg_0_25_41(w_stg_0_25_41, data_operandA[16], data_operandB[25]);
	and stg_0_25_42(w_stg_0_25_42, data_operandA[17], data_operandB[25]);
	and stg_0_25_43(w_stg_0_25_43, data_operandA[18], data_operandB[25]);
	and stg_0_25_44(w_stg_0_25_44, data_operandA[19], data_operandB[25]);
	and stg_0_25_45(w_stg_0_25_45, data_operandA[20], data_operandB[25]);
	and stg_0_25_46(w_stg_0_25_46, data_operandA[21], data_operandB[25]);
	and stg_0_25_47(w_stg_0_25_47, data_operandA[22], data_operandB[25]);
	and stg_0_25_48(w_stg_0_25_48, data_operandA[23], data_operandB[25]);
	and stg_0_25_49(w_stg_0_25_49, data_operandA[24], data_operandB[25]);
	and stg_0_25_50(w_stg_0_25_50, data_operandA[25], data_operandB[25]);
	and stg_0_25_51(w_stg_0_25_51, data_operandA[26], data_operandB[25]);
	and stg_0_25_52(w_stg_0_25_52, data_operandA[27], data_operandB[25]);
	and stg_0_25_53(w_stg_0_25_53, data_operandA[28], data_operandB[25]);
	and stg_0_25_54(w_stg_0_25_54, data_operandA[29], data_operandB[25]);
	and stg_0_25_55(w_stg_0_25_55, data_operandA[30], data_operandB[25]);
	and stg_0_25_56(w_stg_0_25_56, data_operandA[31], data_operandB[25]);
	and stg_0_26_26(w_stg_0_26_26, data_operandA[0], data_operandB[26]);
	and stg_0_26_27(w_stg_0_26_27, data_operandA[1], data_operandB[26]);
	and stg_0_26_28(w_stg_0_26_28, data_operandA[2], data_operandB[26]);
	and stg_0_26_29(w_stg_0_26_29, data_operandA[3], data_operandB[26]);
	and stg_0_26_30(w_stg_0_26_30, data_operandA[4], data_operandB[26]);
	and stg_0_26_31(w_stg_0_26_31, data_operandA[5], data_operandB[26]);
	and stg_0_26_32(w_stg_0_26_32, data_operandA[6], data_operandB[26]);
	and stg_0_26_33(w_stg_0_26_33, data_operandA[7], data_operandB[26]);
	and stg_0_26_34(w_stg_0_26_34, data_operandA[8], data_operandB[26]);
	and stg_0_26_35(w_stg_0_26_35, data_operandA[9], data_operandB[26]);
	and stg_0_26_36(w_stg_0_26_36, data_operandA[10], data_operandB[26]);
	and stg_0_26_37(w_stg_0_26_37, data_operandA[11], data_operandB[26]);
	and stg_0_26_38(w_stg_0_26_38, data_operandA[12], data_operandB[26]);
	and stg_0_26_39(w_stg_0_26_39, data_operandA[13], data_operandB[26]);
	and stg_0_26_40(w_stg_0_26_40, data_operandA[14], data_operandB[26]);
	and stg_0_26_41(w_stg_0_26_41, data_operandA[15], data_operandB[26]);
	and stg_0_26_42(w_stg_0_26_42, data_operandA[16], data_operandB[26]);
	and stg_0_26_43(w_stg_0_26_43, data_operandA[17], data_operandB[26]);
	and stg_0_26_44(w_stg_0_26_44, data_operandA[18], data_operandB[26]);
	and stg_0_26_45(w_stg_0_26_45, data_operandA[19], data_operandB[26]);
	and stg_0_26_46(w_stg_0_26_46, data_operandA[20], data_operandB[26]);
	and stg_0_26_47(w_stg_0_26_47, data_operandA[21], data_operandB[26]);
	and stg_0_26_48(w_stg_0_26_48, data_operandA[22], data_operandB[26]);
	and stg_0_26_49(w_stg_0_26_49, data_operandA[23], data_operandB[26]);
	and stg_0_26_50(w_stg_0_26_50, data_operandA[24], data_operandB[26]);
	and stg_0_26_51(w_stg_0_26_51, data_operandA[25], data_operandB[26]);
	and stg_0_26_52(w_stg_0_26_52, data_operandA[26], data_operandB[26]);
	and stg_0_26_53(w_stg_0_26_53, data_operandA[27], data_operandB[26]);
	and stg_0_26_54(w_stg_0_26_54, data_operandA[28], data_operandB[26]);
	and stg_0_26_55(w_stg_0_26_55, data_operandA[29], data_operandB[26]);
	and stg_0_26_56(w_stg_0_26_56, data_operandA[30], data_operandB[26]);
	and stg_0_26_57(w_stg_0_26_57, data_operandA[31], data_operandB[26]);
	and stg_0_27_27(w_stg_0_27_27, data_operandA[0], data_operandB[27]);
	and stg_0_27_28(w_stg_0_27_28, data_operandA[1], data_operandB[27]);
	and stg_0_27_29(w_stg_0_27_29, data_operandA[2], data_operandB[27]);
	and stg_0_27_30(w_stg_0_27_30, data_operandA[3], data_operandB[27]);
	and stg_0_27_31(w_stg_0_27_31, data_operandA[4], data_operandB[27]);
	and stg_0_27_32(w_stg_0_27_32, data_operandA[5], data_operandB[27]);
	and stg_0_27_33(w_stg_0_27_33, data_operandA[6], data_operandB[27]);
	and stg_0_27_34(w_stg_0_27_34, data_operandA[7], data_operandB[27]);
	and stg_0_27_35(w_stg_0_27_35, data_operandA[8], data_operandB[27]);
	and stg_0_27_36(w_stg_0_27_36, data_operandA[9], data_operandB[27]);
	and stg_0_27_37(w_stg_0_27_37, data_operandA[10], data_operandB[27]);
	and stg_0_27_38(w_stg_0_27_38, data_operandA[11], data_operandB[27]);
	and stg_0_27_39(w_stg_0_27_39, data_operandA[12], data_operandB[27]);
	and stg_0_27_40(w_stg_0_27_40, data_operandA[13], data_operandB[27]);
	and stg_0_27_41(w_stg_0_27_41, data_operandA[14], data_operandB[27]);
	and stg_0_27_42(w_stg_0_27_42, data_operandA[15], data_operandB[27]);
	and stg_0_27_43(w_stg_0_27_43, data_operandA[16], data_operandB[27]);
	and stg_0_27_44(w_stg_0_27_44, data_operandA[17], data_operandB[27]);
	and stg_0_27_45(w_stg_0_27_45, data_operandA[18], data_operandB[27]);
	and stg_0_27_46(w_stg_0_27_46, data_operandA[19], data_operandB[27]);
	and stg_0_27_47(w_stg_0_27_47, data_operandA[20], data_operandB[27]);
	and stg_0_27_48(w_stg_0_27_48, data_operandA[21], data_operandB[27]);
	and stg_0_27_49(w_stg_0_27_49, data_operandA[22], data_operandB[27]);
	and stg_0_27_50(w_stg_0_27_50, data_operandA[23], data_operandB[27]);
	and stg_0_27_51(w_stg_0_27_51, data_operandA[24], data_operandB[27]);
	and stg_0_27_52(w_stg_0_27_52, data_operandA[25], data_operandB[27]);
	and stg_0_27_53(w_stg_0_27_53, data_operandA[26], data_operandB[27]);
	and stg_0_27_54(w_stg_0_27_54, data_operandA[27], data_operandB[27]);
	and stg_0_27_55(w_stg_0_27_55, data_operandA[28], data_operandB[27]);
	and stg_0_27_56(w_stg_0_27_56, data_operandA[29], data_operandB[27]);
	and stg_0_27_57(w_stg_0_27_57, data_operandA[30], data_operandB[27]);
	and stg_0_27_58(w_stg_0_27_58, data_operandA[31], data_operandB[27]);
	and stg_0_28_28(w_stg_0_28_28, data_operandA[0], data_operandB[28]);
	and stg_0_28_29(w_stg_0_28_29, data_operandA[1], data_operandB[28]);
	and stg_0_28_30(w_stg_0_28_30, data_operandA[2], data_operandB[28]);
	and stg_0_28_31(w_stg_0_28_31, data_operandA[3], data_operandB[28]);
	and stg_0_28_32(w_stg_0_28_32, data_operandA[4], data_operandB[28]);
	and stg_0_28_33(w_stg_0_28_33, data_operandA[5], data_operandB[28]);
	and stg_0_28_34(w_stg_0_28_34, data_operandA[6], data_operandB[28]);
	and stg_0_28_35(w_stg_0_28_35, data_operandA[7], data_operandB[28]);
	and stg_0_28_36(w_stg_0_28_36, data_operandA[8], data_operandB[28]);
	and stg_0_28_37(w_stg_0_28_37, data_operandA[9], data_operandB[28]);
	and stg_0_28_38(w_stg_0_28_38, data_operandA[10], data_operandB[28]);
	and stg_0_28_39(w_stg_0_28_39, data_operandA[11], data_operandB[28]);
	and stg_0_28_40(w_stg_0_28_40, data_operandA[12], data_operandB[28]);
	and stg_0_28_41(w_stg_0_28_41, data_operandA[13], data_operandB[28]);
	and stg_0_28_42(w_stg_0_28_42, data_operandA[14], data_operandB[28]);
	and stg_0_28_43(w_stg_0_28_43, data_operandA[15], data_operandB[28]);
	and stg_0_28_44(w_stg_0_28_44, data_operandA[16], data_operandB[28]);
	and stg_0_28_45(w_stg_0_28_45, data_operandA[17], data_operandB[28]);
	and stg_0_28_46(w_stg_0_28_46, data_operandA[18], data_operandB[28]);
	and stg_0_28_47(w_stg_0_28_47, data_operandA[19], data_operandB[28]);
	and stg_0_28_48(w_stg_0_28_48, data_operandA[20], data_operandB[28]);
	and stg_0_28_49(w_stg_0_28_49, data_operandA[21], data_operandB[28]);
	and stg_0_28_50(w_stg_0_28_50, data_operandA[22], data_operandB[28]);
	and stg_0_28_51(w_stg_0_28_51, data_operandA[23], data_operandB[28]);
	and stg_0_28_52(w_stg_0_28_52, data_operandA[24], data_operandB[28]);
	and stg_0_28_53(w_stg_0_28_53, data_operandA[25], data_operandB[28]);
	and stg_0_28_54(w_stg_0_28_54, data_operandA[26], data_operandB[28]);
	and stg_0_28_55(w_stg_0_28_55, data_operandA[27], data_operandB[28]);
	and stg_0_28_56(w_stg_0_28_56, data_operandA[28], data_operandB[28]);
	and stg_0_28_57(w_stg_0_28_57, data_operandA[29], data_operandB[28]);
	and stg_0_28_58(w_stg_0_28_58, data_operandA[30], data_operandB[28]);
	and stg_0_28_59(w_stg_0_28_59, data_operandA[31], data_operandB[28]);
	and stg_0_29_29(w_stg_0_29_29, data_operandA[0], data_operandB[29]);
	and stg_0_29_30(w_stg_0_29_30, data_operandA[1], data_operandB[29]);
	and stg_0_29_31(w_stg_0_29_31, data_operandA[2], data_operandB[29]);
	and stg_0_29_32(w_stg_0_29_32, data_operandA[3], data_operandB[29]);
	and stg_0_29_33(w_stg_0_29_33, data_operandA[4], data_operandB[29]);
	and stg_0_29_34(w_stg_0_29_34, data_operandA[5], data_operandB[29]);
	and stg_0_29_35(w_stg_0_29_35, data_operandA[6], data_operandB[29]);
	and stg_0_29_36(w_stg_0_29_36, data_operandA[7], data_operandB[29]);
	and stg_0_29_37(w_stg_0_29_37, data_operandA[8], data_operandB[29]);
	and stg_0_29_38(w_stg_0_29_38, data_operandA[9], data_operandB[29]);
	and stg_0_29_39(w_stg_0_29_39, data_operandA[10], data_operandB[29]);
	and stg_0_29_40(w_stg_0_29_40, data_operandA[11], data_operandB[29]);
	and stg_0_29_41(w_stg_0_29_41, data_operandA[12], data_operandB[29]);
	and stg_0_29_42(w_stg_0_29_42, data_operandA[13], data_operandB[29]);
	and stg_0_29_43(w_stg_0_29_43, data_operandA[14], data_operandB[29]);
	and stg_0_29_44(w_stg_0_29_44, data_operandA[15], data_operandB[29]);
	and stg_0_29_45(w_stg_0_29_45, data_operandA[16], data_operandB[29]);
	and stg_0_29_46(w_stg_0_29_46, data_operandA[17], data_operandB[29]);
	and stg_0_29_47(w_stg_0_29_47, data_operandA[18], data_operandB[29]);
	and stg_0_29_48(w_stg_0_29_48, data_operandA[19], data_operandB[29]);
	and stg_0_29_49(w_stg_0_29_49, data_operandA[20], data_operandB[29]);
	and stg_0_29_50(w_stg_0_29_50, data_operandA[21], data_operandB[29]);
	and stg_0_29_51(w_stg_0_29_51, data_operandA[22], data_operandB[29]);
	and stg_0_29_52(w_stg_0_29_52, data_operandA[23], data_operandB[29]);
	and stg_0_29_53(w_stg_0_29_53, data_operandA[24], data_operandB[29]);
	and stg_0_29_54(w_stg_0_29_54, data_operandA[25], data_operandB[29]);
	and stg_0_29_55(w_stg_0_29_55, data_operandA[26], data_operandB[29]);
	and stg_0_29_56(w_stg_0_29_56, data_operandA[27], data_operandB[29]);
	and stg_0_29_57(w_stg_0_29_57, data_operandA[28], data_operandB[29]);
	and stg_0_29_58(w_stg_0_29_58, data_operandA[29], data_operandB[29]);
	and stg_0_29_59(w_stg_0_29_59, data_operandA[30], data_operandB[29]);
	and stg_0_29_60(w_stg_0_29_60, data_operandA[31], data_operandB[29]);
	and stg_0_30_30(w_stg_0_30_30, data_operandA[0], data_operandB[30]);
	and stg_0_30_31(w_stg_0_30_31, data_operandA[1], data_operandB[30]);
	and stg_0_30_32(w_stg_0_30_32, data_operandA[2], data_operandB[30]);
	and stg_0_30_33(w_stg_0_30_33, data_operandA[3], data_operandB[30]);
	and stg_0_30_34(w_stg_0_30_34, data_operandA[4], data_operandB[30]);
	and stg_0_30_35(w_stg_0_30_35, data_operandA[5], data_operandB[30]);
	and stg_0_30_36(w_stg_0_30_36, data_operandA[6], data_operandB[30]);
	and stg_0_30_37(w_stg_0_30_37, data_operandA[7], data_operandB[30]);
	and stg_0_30_38(w_stg_0_30_38, data_operandA[8], data_operandB[30]);
	and stg_0_30_39(w_stg_0_30_39, data_operandA[9], data_operandB[30]);
	and stg_0_30_40(w_stg_0_30_40, data_operandA[10], data_operandB[30]);
	and stg_0_30_41(w_stg_0_30_41, data_operandA[11], data_operandB[30]);
	and stg_0_30_42(w_stg_0_30_42, data_operandA[12], data_operandB[30]);
	and stg_0_30_43(w_stg_0_30_43, data_operandA[13], data_operandB[30]);
	and stg_0_30_44(w_stg_0_30_44, data_operandA[14], data_operandB[30]);
	and stg_0_30_45(w_stg_0_30_45, data_operandA[15], data_operandB[30]);
	and stg_0_30_46(w_stg_0_30_46, data_operandA[16], data_operandB[30]);
	and stg_0_30_47(w_stg_0_30_47, data_operandA[17], data_operandB[30]);
	and stg_0_30_48(w_stg_0_30_48, data_operandA[18], data_operandB[30]);
	and stg_0_30_49(w_stg_0_30_49, data_operandA[19], data_operandB[30]);
	and stg_0_30_50(w_stg_0_30_50, data_operandA[20], data_operandB[30]);
	and stg_0_30_51(w_stg_0_30_51, data_operandA[21], data_operandB[30]);
	and stg_0_30_52(w_stg_0_30_52, data_operandA[22], data_operandB[30]);
	and stg_0_30_53(w_stg_0_30_53, data_operandA[23], data_operandB[30]);
	and stg_0_30_54(w_stg_0_30_54, data_operandA[24], data_operandB[30]);
	and stg_0_30_55(w_stg_0_30_55, data_operandA[25], data_operandB[30]);
	and stg_0_30_56(w_stg_0_30_56, data_operandA[26], data_operandB[30]);
	and stg_0_30_57(w_stg_0_30_57, data_operandA[27], data_operandB[30]);
	and stg_0_30_58(w_stg_0_30_58, data_operandA[28], data_operandB[30]);
	and stg_0_30_59(w_stg_0_30_59, data_operandA[29], data_operandB[30]);
	and stg_0_30_60(w_stg_0_30_60, data_operandA[30], data_operandB[30]);
	and stg_0_30_61(w_stg_0_30_61, data_operandA[31], data_operandB[30]);
	and stg_0_31_31(w_stg_0_31_31, data_operandA[0], data_operandB[31]);
	and stg_0_31_32(w_stg_0_31_32, data_operandA[1], data_operandB[31]);
	and stg_0_31_33(w_stg_0_31_33, data_operandA[2], data_operandB[31]);
	and stg_0_31_34(w_stg_0_31_34, data_operandA[3], data_operandB[31]);
	and stg_0_31_35(w_stg_0_31_35, data_operandA[4], data_operandB[31]);
	and stg_0_31_36(w_stg_0_31_36, data_operandA[5], data_operandB[31]);
	and stg_0_31_37(w_stg_0_31_37, data_operandA[6], data_operandB[31]);
	and stg_0_31_38(w_stg_0_31_38, data_operandA[7], data_operandB[31]);
	and stg_0_31_39(w_stg_0_31_39, data_operandA[8], data_operandB[31]);
	and stg_0_31_40(w_stg_0_31_40, data_operandA[9], data_operandB[31]);
	and stg_0_31_41(w_stg_0_31_41, data_operandA[10], data_operandB[31]);
	and stg_0_31_42(w_stg_0_31_42, data_operandA[11], data_operandB[31]);
	and stg_0_31_43(w_stg_0_31_43, data_operandA[12], data_operandB[31]);
	and stg_0_31_44(w_stg_0_31_44, data_operandA[13], data_operandB[31]);
	and stg_0_31_45(w_stg_0_31_45, data_operandA[14], data_operandB[31]);
	and stg_0_31_46(w_stg_0_31_46, data_operandA[15], data_operandB[31]);
	and stg_0_31_47(w_stg_0_31_47, data_operandA[16], data_operandB[31]);
	and stg_0_31_48(w_stg_0_31_48, data_operandA[17], data_operandB[31]);
	and stg_0_31_49(w_stg_0_31_49, data_operandA[18], data_operandB[31]);
	and stg_0_31_50(w_stg_0_31_50, data_operandA[19], data_operandB[31]);
	and stg_0_31_51(w_stg_0_31_51, data_operandA[20], data_operandB[31]);
	and stg_0_31_52(w_stg_0_31_52, data_operandA[21], data_operandB[31]);
	and stg_0_31_53(w_stg_0_31_53, data_operandA[22], data_operandB[31]);
	and stg_0_31_54(w_stg_0_31_54, data_operandA[23], data_operandB[31]);
	and stg_0_31_55(w_stg_0_31_55, data_operandA[24], data_operandB[31]);
	and stg_0_31_56(w_stg_0_31_56, data_operandA[25], data_operandB[31]);
	and stg_0_31_57(w_stg_0_31_57, data_operandA[26], data_operandB[31]);
	and stg_0_31_58(w_stg_0_31_58, data_operandA[27], data_operandB[31]);
	and stg_0_31_59(w_stg_0_31_59, data_operandA[28], data_operandB[31]);
	and stg_0_31_60(w_stg_0_31_60, data_operandA[29], data_operandB[31]);
	and stg_0_31_61(w_stg_0_31_61, data_operandA[30], data_operandB[31]);
	and stg_0_31_62(w_stg_0_31_62, data_operandA[31], data_operandB[31]);
	assign w_stg_1_0_0 = w_stg_0_0_0;
	half_adder ha1( w_stg_1_0_1, w_stg_1_0_2, w_stg_0_0_1, w_stg_0_1_1);
	full_adder_md fa1( w_stg_1_1_2, w_stg_1_0_3, w_stg_0_0_2, w_stg_0_1_2, w_stg_0_2_2);
	full_adder_md fa2( w_stg_1_1_3, w_stg_1_0_4, w_stg_0_0_3, w_stg_0_1_3, w_stg_0_2_3);
	assign w_stg_1_2_3 = w_stg_0_3_3;
	full_adder_md fa3( w_stg_1_1_4, w_stg_1_0_5, w_stg_0_0_4, w_stg_0_1_4, w_stg_0_2_4);
	half_adder ha2( w_stg_1_2_4, w_stg_1_1_5, w_stg_0_3_4, w_stg_0_4_4);
	full_adder_md fa4( w_stg_1_2_5, w_stg_1_0_6, w_stg_0_0_5, w_stg_0_1_5, w_stg_0_2_5);
	full_adder_md fa5( w_stg_1_3_5, w_stg_1_1_6, w_stg_0_3_5, w_stg_0_4_5, w_stg_0_5_5);
	full_adder_md fa6( w_stg_1_2_6, w_stg_1_0_7, w_stg_0_0_6, w_stg_0_1_6, w_stg_0_2_6);
	full_adder_md fa7( w_stg_1_3_6, w_stg_1_1_7, w_stg_0_3_6, w_stg_0_4_6, w_stg_0_5_6);
	assign w_stg_1_4_6 = w_stg_0_6_6;
	full_adder_md fa8( w_stg_1_2_7, w_stg_1_0_8, w_stg_0_0_7, w_stg_0_1_7, w_stg_0_2_7);
	full_adder_md fa9( w_stg_1_3_7, w_stg_1_1_8, w_stg_0_3_7, w_stg_0_4_7, w_stg_0_5_7);
	half_adder ha3( w_stg_1_4_7, w_stg_1_2_8, w_stg_0_6_7, w_stg_0_7_7);
	full_adder_md fa10( w_stg_1_3_8, w_stg_1_0_9, w_stg_0_0_8, w_stg_0_1_8, w_stg_0_2_8);
	full_adder_md fa11( w_stg_1_4_8, w_stg_1_1_9, w_stg_0_3_8, w_stg_0_4_8, w_stg_0_5_8);
	full_adder_md fa12( w_stg_1_5_8, w_stg_1_2_9, w_stg_0_6_8, w_stg_0_7_8, w_stg_0_8_8);
	full_adder_md fa13( w_stg_1_3_9, w_stg_1_0_10, w_stg_0_0_9, w_stg_0_1_9, w_stg_0_2_9);
	full_adder_md fa14( w_stg_1_4_9, w_stg_1_1_10, w_stg_0_3_9, w_stg_0_4_9, w_stg_0_5_9);
	full_adder_md fa15( w_stg_1_5_9, w_stg_1_2_10, w_stg_0_6_9, w_stg_0_7_9, w_stg_0_8_9);
	assign w_stg_1_6_9 = w_stg_0_9_9;
	full_adder_md fa16( w_stg_1_3_10, w_stg_1_0_11, w_stg_0_0_10, w_stg_0_1_10, w_stg_0_2_10);
	full_adder_md fa17( w_stg_1_4_10, w_stg_1_1_11, w_stg_0_3_10, w_stg_0_4_10, w_stg_0_5_10);
	full_adder_md fa18( w_stg_1_5_10, w_stg_1_2_11, w_stg_0_6_10, w_stg_0_7_10, w_stg_0_8_10);
	half_adder ha4( w_stg_1_6_10, w_stg_1_3_11, w_stg_0_9_10, w_stg_0_10_10);
	full_adder_md fa19( w_stg_1_4_11, w_stg_1_0_12, w_stg_0_0_11, w_stg_0_1_11, w_stg_0_2_11);
	full_adder_md fa20( w_stg_1_5_11, w_stg_1_1_12, w_stg_0_3_11, w_stg_0_4_11, w_stg_0_5_11);
	full_adder_md fa21( w_stg_1_6_11, w_stg_1_2_12, w_stg_0_6_11, w_stg_0_7_11, w_stg_0_8_11);
	full_adder_md fa22( w_stg_1_7_11, w_stg_1_3_12, w_stg_0_9_11, w_stg_0_10_11, w_stg_0_11_11);
	full_adder_md fa23( w_stg_1_4_12, w_stg_1_0_13, w_stg_0_0_12, w_stg_0_1_12, w_stg_0_2_12);
	full_adder_md fa24( w_stg_1_5_12, w_stg_1_1_13, w_stg_0_3_12, w_stg_0_4_12, w_stg_0_5_12);
	full_adder_md fa25( w_stg_1_6_12, w_stg_1_2_13, w_stg_0_6_12, w_stg_0_7_12, w_stg_0_8_12);
	full_adder_md fa26( w_stg_1_7_12, w_stg_1_3_13, w_stg_0_9_12, w_stg_0_10_12, w_stg_0_11_12);
	assign w_stg_1_8_12 = w_stg_0_12_12;
	full_adder_md fa27( w_stg_1_4_13, w_stg_1_0_14, w_stg_0_0_13, w_stg_0_1_13, w_stg_0_2_13);
	full_adder_md fa28( w_stg_1_5_13, w_stg_1_1_14, w_stg_0_3_13, w_stg_0_4_13, w_stg_0_5_13);
	full_adder_md fa29( w_stg_1_6_13, w_stg_1_2_14, w_stg_0_6_13, w_stg_0_7_13, w_stg_0_8_13);
	full_adder_md fa30( w_stg_1_7_13, w_stg_1_3_14, w_stg_0_9_13, w_stg_0_10_13, w_stg_0_11_13);
	half_adder ha5( w_stg_1_8_13, w_stg_1_4_14, w_stg_0_12_13, w_stg_0_13_13);
	full_adder_md fa31( w_stg_1_5_14, w_stg_1_0_15, w_stg_0_0_14, w_stg_0_1_14, w_stg_0_2_14);
	full_adder_md fa32( w_stg_1_6_14, w_stg_1_1_15, w_stg_0_3_14, w_stg_0_4_14, w_stg_0_5_14);
	full_adder_md fa33( w_stg_1_7_14, w_stg_1_2_15, w_stg_0_6_14, w_stg_0_7_14, w_stg_0_8_14);
	full_adder_md fa34( w_stg_1_8_14, w_stg_1_3_15, w_stg_0_9_14, w_stg_0_10_14, w_stg_0_11_14);
	full_adder_md fa35( w_stg_1_9_14, w_stg_1_4_15, w_stg_0_12_14, w_stg_0_13_14, w_stg_0_14_14);
	full_adder_md fa36( w_stg_1_5_15, w_stg_1_0_16, w_stg_0_0_15, w_stg_0_1_15, w_stg_0_2_15);
	full_adder_md fa37( w_stg_1_6_15, w_stg_1_1_16, w_stg_0_3_15, w_stg_0_4_15, w_stg_0_5_15);
	full_adder_md fa38( w_stg_1_7_15, w_stg_1_2_16, w_stg_0_6_15, w_stg_0_7_15, w_stg_0_8_15);
	full_adder_md fa39( w_stg_1_8_15, w_stg_1_3_16, w_stg_0_9_15, w_stg_0_10_15, w_stg_0_11_15);
	full_adder_md fa40( w_stg_1_9_15, w_stg_1_4_16, w_stg_0_12_15, w_stg_0_13_15, w_stg_0_14_15);
	assign w_stg_1_10_15 = w_stg_0_15_15;
	full_adder_md fa41( w_stg_1_5_16, w_stg_1_0_17, w_stg_0_0_16, w_stg_0_1_16, w_stg_0_2_16);
	full_adder_md fa42( w_stg_1_6_16, w_stg_1_1_17, w_stg_0_3_16, w_stg_0_4_16, w_stg_0_5_16);
	full_adder_md fa43( w_stg_1_7_16, w_stg_1_2_17, w_stg_0_6_16, w_stg_0_7_16, w_stg_0_8_16);
	full_adder_md fa44( w_stg_1_8_16, w_stg_1_3_17, w_stg_0_9_16, w_stg_0_10_16, w_stg_0_11_16);
	full_adder_md fa45( w_stg_1_9_16, w_stg_1_4_17, w_stg_0_12_16, w_stg_0_13_16, w_stg_0_14_16);
	half_adder ha6( w_stg_1_10_16, w_stg_1_5_17, w_stg_0_15_16, w_stg_0_16_16);
	full_adder_md fa46( w_stg_1_6_17, w_stg_1_0_18, w_stg_0_0_17, w_stg_0_1_17, w_stg_0_2_17);
	full_adder_md fa47( w_stg_1_7_17, w_stg_1_1_18, w_stg_0_3_17, w_stg_0_4_17, w_stg_0_5_17);
	full_adder_md fa48( w_stg_1_8_17, w_stg_1_2_18, w_stg_0_6_17, w_stg_0_7_17, w_stg_0_8_17);
	full_adder_md fa49( w_stg_1_9_17, w_stg_1_3_18, w_stg_0_9_17, w_stg_0_10_17, w_stg_0_11_17);
	full_adder_md fa50( w_stg_1_10_17, w_stg_1_4_18, w_stg_0_12_17, w_stg_0_13_17, w_stg_0_14_17);
	full_adder_md fa51( w_stg_1_11_17, w_stg_1_5_18, w_stg_0_15_17, w_stg_0_16_17, w_stg_0_17_17);
	full_adder_md fa52( w_stg_1_6_18, w_stg_1_0_19, w_stg_0_0_18, w_stg_0_1_18, w_stg_0_2_18);
	full_adder_md fa53( w_stg_1_7_18, w_stg_1_1_19, w_stg_0_3_18, w_stg_0_4_18, w_stg_0_5_18);
	full_adder_md fa54( w_stg_1_8_18, w_stg_1_2_19, w_stg_0_6_18, w_stg_0_7_18, w_stg_0_8_18);
	full_adder_md fa55( w_stg_1_9_18, w_stg_1_3_19, w_stg_0_9_18, w_stg_0_10_18, w_stg_0_11_18);
	full_adder_md fa56( w_stg_1_10_18, w_stg_1_4_19, w_stg_0_12_18, w_stg_0_13_18, w_stg_0_14_18);
	full_adder_md fa57( w_stg_1_11_18, w_stg_1_5_19, w_stg_0_15_18, w_stg_0_16_18, w_stg_0_17_18);
	assign w_stg_1_12_18 = w_stg_0_18_18;
	full_adder_md fa58( w_stg_1_6_19, w_stg_1_0_20, w_stg_0_0_19, w_stg_0_1_19, w_stg_0_2_19);
	full_adder_md fa59( w_stg_1_7_19, w_stg_1_1_20, w_stg_0_3_19, w_stg_0_4_19, w_stg_0_5_19);
	full_adder_md fa60( w_stg_1_8_19, w_stg_1_2_20, w_stg_0_6_19, w_stg_0_7_19, w_stg_0_8_19);
	full_adder_md fa61( w_stg_1_9_19, w_stg_1_3_20, w_stg_0_9_19, w_stg_0_10_19, w_stg_0_11_19);
	full_adder_md fa62( w_stg_1_10_19, w_stg_1_4_20, w_stg_0_12_19, w_stg_0_13_19, w_stg_0_14_19);
	full_adder_md fa63( w_stg_1_11_19, w_stg_1_5_20, w_stg_0_15_19, w_stg_0_16_19, w_stg_0_17_19);
	half_adder ha7( w_stg_1_12_19, w_stg_1_6_20, w_stg_0_18_19, w_stg_0_19_19);
	full_adder_md fa64( w_stg_1_7_20, w_stg_1_0_21, w_stg_0_0_20, w_stg_0_1_20, w_stg_0_2_20);
	full_adder_md fa65( w_stg_1_8_20, w_stg_1_1_21, w_stg_0_3_20, w_stg_0_4_20, w_stg_0_5_20);
	full_adder_md fa66( w_stg_1_9_20, w_stg_1_2_21, w_stg_0_6_20, w_stg_0_7_20, w_stg_0_8_20);
	full_adder_md fa67( w_stg_1_10_20, w_stg_1_3_21, w_stg_0_9_20, w_stg_0_10_20, w_stg_0_11_20);
	full_adder_md fa68( w_stg_1_11_20, w_stg_1_4_21, w_stg_0_12_20, w_stg_0_13_20, w_stg_0_14_20);
	full_adder_md fa69( w_stg_1_12_20, w_stg_1_5_21, w_stg_0_15_20, w_stg_0_16_20, w_stg_0_17_20);
	full_adder_md fa70( w_stg_1_13_20, w_stg_1_6_21, w_stg_0_18_20, w_stg_0_19_20, w_stg_0_20_20);
	full_adder_md fa71( w_stg_1_7_21, w_stg_1_0_22, w_stg_0_0_21, w_stg_0_1_21, w_stg_0_2_21);
	full_adder_md fa72( w_stg_1_8_21, w_stg_1_1_22, w_stg_0_3_21, w_stg_0_4_21, w_stg_0_5_21);
	full_adder_md fa73( w_stg_1_9_21, w_stg_1_2_22, w_stg_0_6_21, w_stg_0_7_21, w_stg_0_8_21);
	full_adder_md fa74( w_stg_1_10_21, w_stg_1_3_22, w_stg_0_9_21, w_stg_0_10_21, w_stg_0_11_21);
	full_adder_md fa75( w_stg_1_11_21, w_stg_1_4_22, w_stg_0_12_21, w_stg_0_13_21, w_stg_0_14_21);
	full_adder_md fa76( w_stg_1_12_21, w_stg_1_5_22, w_stg_0_15_21, w_stg_0_16_21, w_stg_0_17_21);
	full_adder_md fa77( w_stg_1_13_21, w_stg_1_6_22, w_stg_0_18_21, w_stg_0_19_21, w_stg_0_20_21);
	assign w_stg_1_14_21 = w_stg_0_21_21;
	full_adder_md fa78( w_stg_1_7_22, w_stg_1_0_23, w_stg_0_0_22, w_stg_0_1_22, w_stg_0_2_22);
	full_adder_md fa79( w_stg_1_8_22, w_stg_1_1_23, w_stg_0_3_22, w_stg_0_4_22, w_stg_0_5_22);
	full_adder_md fa80( w_stg_1_9_22, w_stg_1_2_23, w_stg_0_6_22, w_stg_0_7_22, w_stg_0_8_22);
	full_adder_md fa81( w_stg_1_10_22, w_stg_1_3_23, w_stg_0_9_22, w_stg_0_10_22, w_stg_0_11_22);
	full_adder_md fa82( w_stg_1_11_22, w_stg_1_4_23, w_stg_0_12_22, w_stg_0_13_22, w_stg_0_14_22);
	full_adder_md fa83( w_stg_1_12_22, w_stg_1_5_23, w_stg_0_15_22, w_stg_0_16_22, w_stg_0_17_22);
	full_adder_md fa84( w_stg_1_13_22, w_stg_1_6_23, w_stg_0_18_22, w_stg_0_19_22, w_stg_0_20_22);
	half_adder ha8( w_stg_1_14_22, w_stg_1_7_23, w_stg_0_21_22, w_stg_0_22_22);
	full_adder_md fa85( w_stg_1_8_23, w_stg_1_0_24, w_stg_0_0_23, w_stg_0_1_23, w_stg_0_2_23);
	full_adder_md fa86( w_stg_1_9_23, w_stg_1_1_24, w_stg_0_3_23, w_stg_0_4_23, w_stg_0_5_23);
	full_adder_md fa87( w_stg_1_10_23, w_stg_1_2_24, w_stg_0_6_23, w_stg_0_7_23, w_stg_0_8_23);
	full_adder_md fa88( w_stg_1_11_23, w_stg_1_3_24, w_stg_0_9_23, w_stg_0_10_23, w_stg_0_11_23);
	full_adder_md fa89( w_stg_1_12_23, w_stg_1_4_24, w_stg_0_12_23, w_stg_0_13_23, w_stg_0_14_23);
	full_adder_md fa90( w_stg_1_13_23, w_stg_1_5_24, w_stg_0_15_23, w_stg_0_16_23, w_stg_0_17_23);
	full_adder_md fa91( w_stg_1_14_23, w_stg_1_6_24, w_stg_0_18_23, w_stg_0_19_23, w_stg_0_20_23);
	full_adder_md fa92( w_stg_1_15_23, w_stg_1_7_24, w_stg_0_21_23, w_stg_0_22_23, w_stg_0_23_23);
	full_adder_md fa93( w_stg_1_8_24, w_stg_1_0_25, w_stg_0_0_24, w_stg_0_1_24, w_stg_0_2_24);
	full_adder_md fa94( w_stg_1_9_24, w_stg_1_1_25, w_stg_0_3_24, w_stg_0_4_24, w_stg_0_5_24);
	full_adder_md fa95( w_stg_1_10_24, w_stg_1_2_25, w_stg_0_6_24, w_stg_0_7_24, w_stg_0_8_24);
	full_adder_md fa96( w_stg_1_11_24, w_stg_1_3_25, w_stg_0_9_24, w_stg_0_10_24, w_stg_0_11_24);
	full_adder_md fa97( w_stg_1_12_24, w_stg_1_4_25, w_stg_0_12_24, w_stg_0_13_24, w_stg_0_14_24);
	full_adder_md fa98( w_stg_1_13_24, w_stg_1_5_25, w_stg_0_15_24, w_stg_0_16_24, w_stg_0_17_24);
	full_adder_md fa99( w_stg_1_14_24, w_stg_1_6_25, w_stg_0_18_24, w_stg_0_19_24, w_stg_0_20_24);
	full_adder_md fa100( w_stg_1_15_24, w_stg_1_7_25, w_stg_0_21_24, w_stg_0_22_24, w_stg_0_23_24);
	assign w_stg_1_16_24 = w_stg_0_24_24;
	full_adder_md fa101( w_stg_1_8_25, w_stg_1_0_26, w_stg_0_0_25, w_stg_0_1_25, w_stg_0_2_25);
	full_adder_md fa102( w_stg_1_9_25, w_stg_1_1_26, w_stg_0_3_25, w_stg_0_4_25, w_stg_0_5_25);
	full_adder_md fa103( w_stg_1_10_25, w_stg_1_2_26, w_stg_0_6_25, w_stg_0_7_25, w_stg_0_8_25);
	full_adder_md fa104( w_stg_1_11_25, w_stg_1_3_26, w_stg_0_9_25, w_stg_0_10_25, w_stg_0_11_25);
	full_adder_md fa105( w_stg_1_12_25, w_stg_1_4_26, w_stg_0_12_25, w_stg_0_13_25, w_stg_0_14_25);
	full_adder_md fa106( w_stg_1_13_25, w_stg_1_5_26, w_stg_0_15_25, w_stg_0_16_25, w_stg_0_17_25);
	full_adder_md fa107( w_stg_1_14_25, w_stg_1_6_26, w_stg_0_18_25, w_stg_0_19_25, w_stg_0_20_25);
	full_adder_md fa108( w_stg_1_15_25, w_stg_1_7_26, w_stg_0_21_25, w_stg_0_22_25, w_stg_0_23_25);
	half_adder ha9( w_stg_1_16_25, w_stg_1_8_26, w_stg_0_24_25, w_stg_0_25_25);
	full_adder_md fa109( w_stg_1_9_26, w_stg_1_0_27, w_stg_0_0_26, w_stg_0_1_26, w_stg_0_2_26);
	full_adder_md fa110( w_stg_1_10_26, w_stg_1_1_27, w_stg_0_3_26, w_stg_0_4_26, w_stg_0_5_26);
	full_adder_md fa111( w_stg_1_11_26, w_stg_1_2_27, w_stg_0_6_26, w_stg_0_7_26, w_stg_0_8_26);
	full_adder_md fa112( w_stg_1_12_26, w_stg_1_3_27, w_stg_0_9_26, w_stg_0_10_26, w_stg_0_11_26);
	full_adder_md fa113( w_stg_1_13_26, w_stg_1_4_27, w_stg_0_12_26, w_stg_0_13_26, w_stg_0_14_26);
	full_adder_md fa114( w_stg_1_14_26, w_stg_1_5_27, w_stg_0_15_26, w_stg_0_16_26, w_stg_0_17_26);
	full_adder_md fa115( w_stg_1_15_26, w_stg_1_6_27, w_stg_0_18_26, w_stg_0_19_26, w_stg_0_20_26);
	full_adder_md fa116( w_stg_1_16_26, w_stg_1_7_27, w_stg_0_21_26, w_stg_0_22_26, w_stg_0_23_26);
	full_adder_md fa117( w_stg_1_17_26, w_stg_1_8_27, w_stg_0_24_26, w_stg_0_25_26, w_stg_0_26_26);
	full_adder_md fa118( w_stg_1_9_27, w_stg_1_0_28, w_stg_0_0_27, w_stg_0_1_27, w_stg_0_2_27);
	full_adder_md fa119( w_stg_1_10_27, w_stg_1_1_28, w_stg_0_3_27, w_stg_0_4_27, w_stg_0_5_27);
	full_adder_md fa120( w_stg_1_11_27, w_stg_1_2_28, w_stg_0_6_27, w_stg_0_7_27, w_stg_0_8_27);
	full_adder_md fa121( w_stg_1_12_27, w_stg_1_3_28, w_stg_0_9_27, w_stg_0_10_27, w_stg_0_11_27);
	full_adder_md fa122( w_stg_1_13_27, w_stg_1_4_28, w_stg_0_12_27, w_stg_0_13_27, w_stg_0_14_27);
	full_adder_md fa123( w_stg_1_14_27, w_stg_1_5_28, w_stg_0_15_27, w_stg_0_16_27, w_stg_0_17_27);
	full_adder_md fa124( w_stg_1_15_27, w_stg_1_6_28, w_stg_0_18_27, w_stg_0_19_27, w_stg_0_20_27);
	full_adder_md fa125( w_stg_1_16_27, w_stg_1_7_28, w_stg_0_21_27, w_stg_0_22_27, w_stg_0_23_27);
	full_adder_md fa126( w_stg_1_17_27, w_stg_1_8_28, w_stg_0_24_27, w_stg_0_25_27, w_stg_0_26_27);
	assign w_stg_1_18_27 = w_stg_0_27_27;
	full_adder_md fa127( w_stg_1_9_28, w_stg_1_0_29, w_stg_0_0_28, w_stg_0_1_28, w_stg_0_2_28);
	full_adder_md fa128( w_stg_1_10_28, w_stg_1_1_29, w_stg_0_3_28, w_stg_0_4_28, w_stg_0_5_28);
	full_adder_md fa129( w_stg_1_11_28, w_stg_1_2_29, w_stg_0_6_28, w_stg_0_7_28, w_stg_0_8_28);
	full_adder_md fa130( w_stg_1_12_28, w_stg_1_3_29, w_stg_0_9_28, w_stg_0_10_28, w_stg_0_11_28);
	full_adder_md fa131( w_stg_1_13_28, w_stg_1_4_29, w_stg_0_12_28, w_stg_0_13_28, w_stg_0_14_28);
	full_adder_md fa132( w_stg_1_14_28, w_stg_1_5_29, w_stg_0_15_28, w_stg_0_16_28, w_stg_0_17_28);
	full_adder_md fa133( w_stg_1_15_28, w_stg_1_6_29, w_stg_0_18_28, w_stg_0_19_28, w_stg_0_20_28);
	full_adder_md fa134( w_stg_1_16_28, w_stg_1_7_29, w_stg_0_21_28, w_stg_0_22_28, w_stg_0_23_28);
	full_adder_md fa135( w_stg_1_17_28, w_stg_1_8_29, w_stg_0_24_28, w_stg_0_25_28, w_stg_0_26_28);
	half_adder ha10( w_stg_1_18_28, w_stg_1_9_29, w_stg_0_27_28, w_stg_0_28_28);
	full_adder_md fa136( w_stg_1_10_29, w_stg_1_0_30, w_stg_0_0_29, w_stg_0_1_29, w_stg_0_2_29);
	full_adder_md fa137( w_stg_1_11_29, w_stg_1_1_30, w_stg_0_3_29, w_stg_0_4_29, w_stg_0_5_29);
	full_adder_md fa138( w_stg_1_12_29, w_stg_1_2_30, w_stg_0_6_29, w_stg_0_7_29, w_stg_0_8_29);
	full_adder_md fa139( w_stg_1_13_29, w_stg_1_3_30, w_stg_0_9_29, w_stg_0_10_29, w_stg_0_11_29);
	full_adder_md fa140( w_stg_1_14_29, w_stg_1_4_30, w_stg_0_12_29, w_stg_0_13_29, w_stg_0_14_29);
	full_adder_md fa141( w_stg_1_15_29, w_stg_1_5_30, w_stg_0_15_29, w_stg_0_16_29, w_stg_0_17_29);
	full_adder_md fa142( w_stg_1_16_29, w_stg_1_6_30, w_stg_0_18_29, w_stg_0_19_29, w_stg_0_20_29);
	full_adder_md fa143( w_stg_1_17_29, w_stg_1_7_30, w_stg_0_21_29, w_stg_0_22_29, w_stg_0_23_29);
	full_adder_md fa144( w_stg_1_18_29, w_stg_1_8_30, w_stg_0_24_29, w_stg_0_25_29, w_stg_0_26_29);
	full_adder_md fa145( w_stg_1_19_29, w_stg_1_9_30, w_stg_0_27_29, w_stg_0_28_29, w_stg_0_29_29);
	full_adder_md fa146( w_stg_1_10_30, w_stg_1_0_31, w_stg_0_0_30, w_stg_0_1_30, w_stg_0_2_30);
	full_adder_md fa147( w_stg_1_11_30, w_stg_1_1_31, w_stg_0_3_30, w_stg_0_4_30, w_stg_0_5_30);
	full_adder_md fa148( w_stg_1_12_30, w_stg_1_2_31, w_stg_0_6_30, w_stg_0_7_30, w_stg_0_8_30);
	full_adder_md fa149( w_stg_1_13_30, w_stg_1_3_31, w_stg_0_9_30, w_stg_0_10_30, w_stg_0_11_30);
	full_adder_md fa150( w_stg_1_14_30, w_stg_1_4_31, w_stg_0_12_30, w_stg_0_13_30, w_stg_0_14_30);
	full_adder_md fa151( w_stg_1_15_30, w_stg_1_5_31, w_stg_0_15_30, w_stg_0_16_30, w_stg_0_17_30);
	full_adder_md fa152( w_stg_1_16_30, w_stg_1_6_31, w_stg_0_18_30, w_stg_0_19_30, w_stg_0_20_30);
	full_adder_md fa153( w_stg_1_17_30, w_stg_1_7_31, w_stg_0_21_30, w_stg_0_22_30, w_stg_0_23_30);
	full_adder_md fa154( w_stg_1_18_30, w_stg_1_8_31, w_stg_0_24_30, w_stg_0_25_30, w_stg_0_26_30);
	full_adder_md fa155( w_stg_1_19_30, w_stg_1_9_31, w_stg_0_27_30, w_stg_0_28_30, w_stg_0_29_30);
	assign w_stg_1_20_30 = w_stg_0_30_30;
	full_adder_md fa156( w_stg_1_10_31, w_stg_1_0_32, w_stg_0_0_31, w_stg_0_1_31, w_stg_0_2_31);
	full_adder_md fa157( w_stg_1_11_31, w_stg_1_1_32, w_stg_0_3_31, w_stg_0_4_31, w_stg_0_5_31);
	full_adder_md fa158( w_stg_1_12_31, w_stg_1_2_32, w_stg_0_6_31, w_stg_0_7_31, w_stg_0_8_31);
	full_adder_md fa159( w_stg_1_13_31, w_stg_1_3_32, w_stg_0_9_31, w_stg_0_10_31, w_stg_0_11_31);
	full_adder_md fa160( w_stg_1_14_31, w_stg_1_4_32, w_stg_0_12_31, w_stg_0_13_31, w_stg_0_14_31);
	full_adder_md fa161( w_stg_1_15_31, w_stg_1_5_32, w_stg_0_15_31, w_stg_0_16_31, w_stg_0_17_31);
	full_adder_md fa162( w_stg_1_16_31, w_stg_1_6_32, w_stg_0_18_31, w_stg_0_19_31, w_stg_0_20_31);
	full_adder_md fa163( w_stg_1_17_31, w_stg_1_7_32, w_stg_0_21_31, w_stg_0_22_31, w_stg_0_23_31);
	full_adder_md fa164( w_stg_1_18_31, w_stg_1_8_32, w_stg_0_24_31, w_stg_0_25_31, w_stg_0_26_31);
	full_adder_md fa165( w_stg_1_19_31, w_stg_1_9_32, w_stg_0_27_31, w_stg_0_28_31, w_stg_0_29_31);
	half_adder ha11( w_stg_1_20_31, w_stg_1_10_32, w_stg_0_30_31, w_stg_0_31_31);
	half_adder ha12( w_stg_1_11_32, w_stg_1_0_33, w_stg_0_1_32, w_stg_0_2_32);
	full_adder_md fa166( w_stg_1_12_32, w_stg_1_1_33, w_stg_0_3_32, w_stg_0_4_32, w_stg_0_5_32);
	full_adder_md fa167( w_stg_1_13_32, w_stg_1_2_33, w_stg_0_6_32, w_stg_0_7_32, w_stg_0_8_32);
	full_adder_md fa168( w_stg_1_14_32, w_stg_1_3_33, w_stg_0_9_32, w_stg_0_10_32, w_stg_0_11_32);
	full_adder_md fa169( w_stg_1_15_32, w_stg_1_4_33, w_stg_0_12_32, w_stg_0_13_32, w_stg_0_14_32);
	full_adder_md fa170( w_stg_1_16_32, w_stg_1_5_33, w_stg_0_15_32, w_stg_0_16_32, w_stg_0_17_32);
	full_adder_md fa171( w_stg_1_17_32, w_stg_1_6_33, w_stg_0_18_32, w_stg_0_19_32, w_stg_0_20_32);
	full_adder_md fa172( w_stg_1_18_32, w_stg_1_7_33, w_stg_0_21_32, w_stg_0_22_32, w_stg_0_23_32);
	full_adder_md fa173( w_stg_1_19_32, w_stg_1_8_33, w_stg_0_24_32, w_stg_0_25_32, w_stg_0_26_32);
	full_adder_md fa174( w_stg_1_20_32, w_stg_1_9_33, w_stg_0_27_32, w_stg_0_28_32, w_stg_0_29_32);
	half_adder ha13( w_stg_1_21_32, w_stg_1_10_33, w_stg_0_30_32, w_stg_0_31_32);
	assign w_stg_1_11_33 = w_stg_0_2_33;
	full_adder_md fa175( w_stg_1_12_33, w_stg_1_0_34, w_stg_0_3_33, w_stg_0_4_33, w_stg_0_5_33);
	full_adder_md fa176( w_stg_1_13_33, w_stg_1_1_34, w_stg_0_6_33, w_stg_0_7_33, w_stg_0_8_33);
	full_adder_md fa177( w_stg_1_14_33, w_stg_1_2_34, w_stg_0_9_33, w_stg_0_10_33, w_stg_0_11_33);
	full_adder_md fa178( w_stg_1_15_33, w_stg_1_3_34, w_stg_0_12_33, w_stg_0_13_33, w_stg_0_14_33);
	full_adder_md fa179( w_stg_1_16_33, w_stg_1_4_34, w_stg_0_15_33, w_stg_0_16_33, w_stg_0_17_33);
	full_adder_md fa180( w_stg_1_17_33, w_stg_1_5_34, w_stg_0_18_33, w_stg_0_19_33, w_stg_0_20_33);
	full_adder_md fa181( w_stg_1_18_33, w_stg_1_6_34, w_stg_0_21_33, w_stg_0_22_33, w_stg_0_23_33);
	full_adder_md fa182( w_stg_1_19_33, w_stg_1_7_34, w_stg_0_24_33, w_stg_0_25_33, w_stg_0_26_33);
	full_adder_md fa183( w_stg_1_20_33, w_stg_1_8_34, w_stg_0_27_33, w_stg_0_28_33, w_stg_0_29_33);
	half_adder ha14( w_stg_1_21_33, w_stg_1_9_34, w_stg_0_30_33, w_stg_0_31_33);
	full_adder_md fa184( w_stg_1_10_34, w_stg_1_0_35, w_stg_0_3_34, w_stg_0_4_34, w_stg_0_5_34);
	full_adder_md fa185( w_stg_1_11_34, w_stg_1_1_35, w_stg_0_6_34, w_stg_0_7_34, w_stg_0_8_34);
	full_adder_md fa186( w_stg_1_12_34, w_stg_1_2_35, w_stg_0_9_34, w_stg_0_10_34, w_stg_0_11_34);
	full_adder_md fa187( w_stg_1_13_34, w_stg_1_3_35, w_stg_0_12_34, w_stg_0_13_34, w_stg_0_14_34);
	full_adder_md fa188( w_stg_1_14_34, w_stg_1_4_35, w_stg_0_15_34, w_stg_0_16_34, w_stg_0_17_34);
	full_adder_md fa189( w_stg_1_15_34, w_stg_1_5_35, w_stg_0_18_34, w_stg_0_19_34, w_stg_0_20_34);
	full_adder_md fa190( w_stg_1_16_34, w_stg_1_6_35, w_stg_0_21_34, w_stg_0_22_34, w_stg_0_23_34);
	full_adder_md fa191( w_stg_1_17_34, w_stg_1_7_35, w_stg_0_24_34, w_stg_0_25_34, w_stg_0_26_34);
	full_adder_md fa192( w_stg_1_18_34, w_stg_1_8_35, w_stg_0_27_34, w_stg_0_28_34, w_stg_0_29_34);
	half_adder ha15( w_stg_1_19_34, w_stg_1_9_35, w_stg_0_30_34, w_stg_0_31_34);
	half_adder ha16( w_stg_1_10_35, w_stg_1_0_36, w_stg_0_4_35, w_stg_0_5_35);
	full_adder_md fa193( w_stg_1_11_35, w_stg_1_1_36, w_stg_0_6_35, w_stg_0_7_35, w_stg_0_8_35);
	full_adder_md fa194( w_stg_1_12_35, w_stg_1_2_36, w_stg_0_9_35, w_stg_0_10_35, w_stg_0_11_35);
	full_adder_md fa195( w_stg_1_13_35, w_stg_1_3_36, w_stg_0_12_35, w_stg_0_13_35, w_stg_0_14_35);
	full_adder_md fa196( w_stg_1_14_35, w_stg_1_4_36, w_stg_0_15_35, w_stg_0_16_35, w_stg_0_17_35);
	full_adder_md fa197( w_stg_1_15_35, w_stg_1_5_36, w_stg_0_18_35, w_stg_0_19_35, w_stg_0_20_35);
	full_adder_md fa198( w_stg_1_16_35, w_stg_1_6_36, w_stg_0_21_35, w_stg_0_22_35, w_stg_0_23_35);
	full_adder_md fa199( w_stg_1_17_35, w_stg_1_7_36, w_stg_0_24_35, w_stg_0_25_35, w_stg_0_26_35);
	full_adder_md fa200( w_stg_1_18_35, w_stg_1_8_36, w_stg_0_27_35, w_stg_0_28_35, w_stg_0_29_35);
	half_adder ha17( w_stg_1_19_35, w_stg_1_9_36, w_stg_0_30_35, w_stg_0_31_35);
	assign w_stg_1_10_36 = w_stg_0_5_36;
	full_adder_md fa201( w_stg_1_11_36, w_stg_1_0_37, w_stg_0_6_36, w_stg_0_7_36, w_stg_0_8_36);
	full_adder_md fa202( w_stg_1_12_36, w_stg_1_1_37, w_stg_0_9_36, w_stg_0_10_36, w_stg_0_11_36);
	full_adder_md fa203( w_stg_1_13_36, w_stg_1_2_37, w_stg_0_12_36, w_stg_0_13_36, w_stg_0_14_36);
	full_adder_md fa204( w_stg_1_14_36, w_stg_1_3_37, w_stg_0_15_36, w_stg_0_16_36, w_stg_0_17_36);
	full_adder_md fa205( w_stg_1_15_36, w_stg_1_4_37, w_stg_0_18_36, w_stg_0_19_36, w_stg_0_20_36);
	full_adder_md fa206( w_stg_1_16_36, w_stg_1_5_37, w_stg_0_21_36, w_stg_0_22_36, w_stg_0_23_36);
	full_adder_md fa207( w_stg_1_17_36, w_stg_1_6_37, w_stg_0_24_36, w_stg_0_25_36, w_stg_0_26_36);
	full_adder_md fa208( w_stg_1_18_36, w_stg_1_7_37, w_stg_0_27_36, w_stg_0_28_36, w_stg_0_29_36);
	half_adder ha18( w_stg_1_19_36, w_stg_1_8_37, w_stg_0_30_36, w_stg_0_31_36);
	full_adder_md fa209( w_stg_1_9_37, w_stg_1_0_38, w_stg_0_6_37, w_stg_0_7_37, w_stg_0_8_37);
	full_adder_md fa210( w_stg_1_10_37, w_stg_1_1_38, w_stg_0_9_37, w_stg_0_10_37, w_stg_0_11_37);
	full_adder_md fa211( w_stg_1_11_37, w_stg_1_2_38, w_stg_0_12_37, w_stg_0_13_37, w_stg_0_14_37);
	full_adder_md fa212( w_stg_1_12_37, w_stg_1_3_38, w_stg_0_15_37, w_stg_0_16_37, w_stg_0_17_37);
	full_adder_md fa213( w_stg_1_13_37, w_stg_1_4_38, w_stg_0_18_37, w_stg_0_19_37, w_stg_0_20_37);
	full_adder_md fa214( w_stg_1_14_37, w_stg_1_5_38, w_stg_0_21_37, w_stg_0_22_37, w_stg_0_23_37);
	full_adder_md fa215( w_stg_1_15_37, w_stg_1_6_38, w_stg_0_24_37, w_stg_0_25_37, w_stg_0_26_37);
	full_adder_md fa216( w_stg_1_16_37, w_stg_1_7_38, w_stg_0_27_37, w_stg_0_28_37, w_stg_0_29_37);
	half_adder ha19( w_stg_1_17_37, w_stg_1_8_38, w_stg_0_30_37, w_stg_0_31_37);
	half_adder ha20( w_stg_1_9_38, w_stg_1_0_39, w_stg_0_7_38, w_stg_0_8_38);
	full_adder_md fa217( w_stg_1_10_38, w_stg_1_1_39, w_stg_0_9_38, w_stg_0_10_38, w_stg_0_11_38);
	full_adder_md fa218( w_stg_1_11_38, w_stg_1_2_39, w_stg_0_12_38, w_stg_0_13_38, w_stg_0_14_38);
	full_adder_md fa219( w_stg_1_12_38, w_stg_1_3_39, w_stg_0_15_38, w_stg_0_16_38, w_stg_0_17_38);
	full_adder_md fa220( w_stg_1_13_38, w_stg_1_4_39, w_stg_0_18_38, w_stg_0_19_38, w_stg_0_20_38);
	full_adder_md fa221( w_stg_1_14_38, w_stg_1_5_39, w_stg_0_21_38, w_stg_0_22_38, w_stg_0_23_38);
	full_adder_md fa222( w_stg_1_15_38, w_stg_1_6_39, w_stg_0_24_38, w_stg_0_25_38, w_stg_0_26_38);
	full_adder_md fa223( w_stg_1_16_38, w_stg_1_7_39, w_stg_0_27_38, w_stg_0_28_38, w_stg_0_29_38);
	half_adder ha21( w_stg_1_17_38, w_stg_1_8_39, w_stg_0_30_38, w_stg_0_31_38);
	assign w_stg_1_9_39 = w_stg_0_8_39;
	full_adder_md fa224( w_stg_1_10_39, w_stg_1_0_40, w_stg_0_9_39, w_stg_0_10_39, w_stg_0_11_39);
	full_adder_md fa225( w_stg_1_11_39, w_stg_1_1_40, w_stg_0_12_39, w_stg_0_13_39, w_stg_0_14_39);
	full_adder_md fa226( w_stg_1_12_39, w_stg_1_2_40, w_stg_0_15_39, w_stg_0_16_39, w_stg_0_17_39);
	full_adder_md fa227( w_stg_1_13_39, w_stg_1_3_40, w_stg_0_18_39, w_stg_0_19_39, w_stg_0_20_39);
	full_adder_md fa228( w_stg_1_14_39, w_stg_1_4_40, w_stg_0_21_39, w_stg_0_22_39, w_stg_0_23_39);
	full_adder_md fa229( w_stg_1_15_39, w_stg_1_5_40, w_stg_0_24_39, w_stg_0_25_39, w_stg_0_26_39);
	full_adder_md fa230( w_stg_1_16_39, w_stg_1_6_40, w_stg_0_27_39, w_stg_0_28_39, w_stg_0_29_39);
	half_adder ha22( w_stg_1_17_39, w_stg_1_7_40, w_stg_0_30_39, w_stg_0_31_39);
	full_adder_md fa231( w_stg_1_8_40, w_stg_1_0_41, w_stg_0_9_40, w_stg_0_10_40, w_stg_0_11_40);
	full_adder_md fa232( w_stg_1_9_40, w_stg_1_1_41, w_stg_0_12_40, w_stg_0_13_40, w_stg_0_14_40);
	full_adder_md fa233( w_stg_1_10_40, w_stg_1_2_41, w_stg_0_15_40, w_stg_0_16_40, w_stg_0_17_40);
	full_adder_md fa234( w_stg_1_11_40, w_stg_1_3_41, w_stg_0_18_40, w_stg_0_19_40, w_stg_0_20_40);
	full_adder_md fa235( w_stg_1_12_40, w_stg_1_4_41, w_stg_0_21_40, w_stg_0_22_40, w_stg_0_23_40);
	full_adder_md fa236( w_stg_1_13_40, w_stg_1_5_41, w_stg_0_24_40, w_stg_0_25_40, w_stg_0_26_40);
	full_adder_md fa237( w_stg_1_14_40, w_stg_1_6_41, w_stg_0_27_40, w_stg_0_28_40, w_stg_0_29_40);
	half_adder ha23( w_stg_1_15_40, w_stg_1_7_41, w_stg_0_30_40, w_stg_0_31_40);
	half_adder ha24( w_stg_1_8_41, w_stg_1_0_42, w_stg_0_10_41, w_stg_0_11_41);
	full_adder_md fa238( w_stg_1_9_41, w_stg_1_1_42, w_stg_0_12_41, w_stg_0_13_41, w_stg_0_14_41);
	full_adder_md fa239( w_stg_1_10_41, w_stg_1_2_42, w_stg_0_15_41, w_stg_0_16_41, w_stg_0_17_41);
	full_adder_md fa240( w_stg_1_11_41, w_stg_1_3_42, w_stg_0_18_41, w_stg_0_19_41, w_stg_0_20_41);
	full_adder_md fa241( w_stg_1_12_41, w_stg_1_4_42, w_stg_0_21_41, w_stg_0_22_41, w_stg_0_23_41);
	full_adder_md fa242( w_stg_1_13_41, w_stg_1_5_42, w_stg_0_24_41, w_stg_0_25_41, w_stg_0_26_41);
	full_adder_md fa243( w_stg_1_14_41, w_stg_1_6_42, w_stg_0_27_41, w_stg_0_28_41, w_stg_0_29_41);
	half_adder ha25( w_stg_1_15_41, w_stg_1_7_42, w_stg_0_30_41, w_stg_0_31_41);
	assign w_stg_1_8_42 = w_stg_0_11_42;
	full_adder_md fa244( w_stg_1_9_42, w_stg_1_0_43, w_stg_0_12_42, w_stg_0_13_42, w_stg_0_14_42);
	full_adder_md fa245( w_stg_1_10_42, w_stg_1_1_43, w_stg_0_15_42, w_stg_0_16_42, w_stg_0_17_42);
	full_adder_md fa246( w_stg_1_11_42, w_stg_1_2_43, w_stg_0_18_42, w_stg_0_19_42, w_stg_0_20_42);
	full_adder_md fa247( w_stg_1_12_42, w_stg_1_3_43, w_stg_0_21_42, w_stg_0_22_42, w_stg_0_23_42);
	full_adder_md fa248( w_stg_1_13_42, w_stg_1_4_43, w_stg_0_24_42, w_stg_0_25_42, w_stg_0_26_42);
	full_adder_md fa249( w_stg_1_14_42, w_stg_1_5_43, w_stg_0_27_42, w_stg_0_28_42, w_stg_0_29_42);
	half_adder ha26( w_stg_1_15_42, w_stg_1_6_43, w_stg_0_30_42, w_stg_0_31_42);
	full_adder_md fa250( w_stg_1_7_43, w_stg_1_0_44, w_stg_0_12_43, w_stg_0_13_43, w_stg_0_14_43);
	full_adder_md fa251( w_stg_1_8_43, w_stg_1_1_44, w_stg_0_15_43, w_stg_0_16_43, w_stg_0_17_43);
	full_adder_md fa252( w_stg_1_9_43, w_stg_1_2_44, w_stg_0_18_43, w_stg_0_19_43, w_stg_0_20_43);
	full_adder_md fa253( w_stg_1_10_43, w_stg_1_3_44, w_stg_0_21_43, w_stg_0_22_43, w_stg_0_23_43);
	full_adder_md fa254( w_stg_1_11_43, w_stg_1_4_44, w_stg_0_24_43, w_stg_0_25_43, w_stg_0_26_43);
	full_adder_md fa255( w_stg_1_12_43, w_stg_1_5_44, w_stg_0_27_43, w_stg_0_28_43, w_stg_0_29_43);
	half_adder ha27( w_stg_1_13_43, w_stg_1_6_44, w_stg_0_30_43, w_stg_0_31_43);
	half_adder ha28( w_stg_1_7_44, w_stg_1_0_45, w_stg_0_13_44, w_stg_0_14_44);
	full_adder_md fa256( w_stg_1_8_44, w_stg_1_1_45, w_stg_0_15_44, w_stg_0_16_44, w_stg_0_17_44);
	full_adder_md fa257( w_stg_1_9_44, w_stg_1_2_45, w_stg_0_18_44, w_stg_0_19_44, w_stg_0_20_44);
	full_adder_md fa258( w_stg_1_10_44, w_stg_1_3_45, w_stg_0_21_44, w_stg_0_22_44, w_stg_0_23_44);
	full_adder_md fa259( w_stg_1_11_44, w_stg_1_4_45, w_stg_0_24_44, w_stg_0_25_44, w_stg_0_26_44);
	full_adder_md fa260( w_stg_1_12_44, w_stg_1_5_45, w_stg_0_27_44, w_stg_0_28_44, w_stg_0_29_44);
	half_adder ha29( w_stg_1_13_44, w_stg_1_6_45, w_stg_0_30_44, w_stg_0_31_44);
	assign w_stg_1_7_45 = w_stg_0_14_45;
	full_adder_md fa261( w_stg_1_8_45, w_stg_1_0_46, w_stg_0_15_45, w_stg_0_16_45, w_stg_0_17_45);
	full_adder_md fa262( w_stg_1_9_45, w_stg_1_1_46, w_stg_0_18_45, w_stg_0_19_45, w_stg_0_20_45);
	full_adder_md fa263( w_stg_1_10_45, w_stg_1_2_46, w_stg_0_21_45, w_stg_0_22_45, w_stg_0_23_45);
	full_adder_md fa264( w_stg_1_11_45, w_stg_1_3_46, w_stg_0_24_45, w_stg_0_25_45, w_stg_0_26_45);
	full_adder_md fa265( w_stg_1_12_45, w_stg_1_4_46, w_stg_0_27_45, w_stg_0_28_45, w_stg_0_29_45);
	half_adder ha30( w_stg_1_13_45, w_stg_1_5_46, w_stg_0_30_45, w_stg_0_31_45);
	full_adder_md fa266( w_stg_1_6_46, w_stg_1_0_47, w_stg_0_15_46, w_stg_0_16_46, w_stg_0_17_46);
	full_adder_md fa267( w_stg_1_7_46, w_stg_1_1_47, w_stg_0_18_46, w_stg_0_19_46, w_stg_0_20_46);
	full_adder_md fa268( w_stg_1_8_46, w_stg_1_2_47, w_stg_0_21_46, w_stg_0_22_46, w_stg_0_23_46);
	full_adder_md fa269( w_stg_1_9_46, w_stg_1_3_47, w_stg_0_24_46, w_stg_0_25_46, w_stg_0_26_46);
	full_adder_md fa270( w_stg_1_10_46, w_stg_1_4_47, w_stg_0_27_46, w_stg_0_28_46, w_stg_0_29_46);
	half_adder ha31( w_stg_1_11_46, w_stg_1_5_47, w_stg_0_30_46, w_stg_0_31_46);
	half_adder ha32( w_stg_1_6_47, w_stg_1_0_48, w_stg_0_16_47, w_stg_0_17_47);
	full_adder_md fa271( w_stg_1_7_47, w_stg_1_1_48, w_stg_0_18_47, w_stg_0_19_47, w_stg_0_20_47);
	full_adder_md fa272( w_stg_1_8_47, w_stg_1_2_48, w_stg_0_21_47, w_stg_0_22_47, w_stg_0_23_47);
	full_adder_md fa273( w_stg_1_9_47, w_stg_1_3_48, w_stg_0_24_47, w_stg_0_25_47, w_stg_0_26_47);
	full_adder_md fa274( w_stg_1_10_47, w_stg_1_4_48, w_stg_0_27_47, w_stg_0_28_47, w_stg_0_29_47);
	half_adder ha33( w_stg_1_11_47, w_stg_1_5_48, w_stg_0_30_47, w_stg_0_31_47);
	assign w_stg_1_6_48 = w_stg_0_17_48;
	full_adder_md fa275( w_stg_1_7_48, w_stg_1_0_49, w_stg_0_18_48, w_stg_0_19_48, w_stg_0_20_48);
	full_adder_md fa276( w_stg_1_8_48, w_stg_1_1_49, w_stg_0_21_48, w_stg_0_22_48, w_stg_0_23_48);
	full_adder_md fa277( w_stg_1_9_48, w_stg_1_2_49, w_stg_0_24_48, w_stg_0_25_48, w_stg_0_26_48);
	full_adder_md fa278( w_stg_1_10_48, w_stg_1_3_49, w_stg_0_27_48, w_stg_0_28_48, w_stg_0_29_48);
	half_adder ha34( w_stg_1_11_48, w_stg_1_4_49, w_stg_0_30_48, w_stg_0_31_48);
	full_adder_md fa279( w_stg_1_5_49, w_stg_1_0_50, w_stg_0_18_49, w_stg_0_19_49, w_stg_0_20_49);
	full_adder_md fa280( w_stg_1_6_49, w_stg_1_1_50, w_stg_0_21_49, w_stg_0_22_49, w_stg_0_23_49);
	full_adder_md fa281( w_stg_1_7_49, w_stg_1_2_50, w_stg_0_24_49, w_stg_0_25_49, w_stg_0_26_49);
	full_adder_md fa282( w_stg_1_8_49, w_stg_1_3_50, w_stg_0_27_49, w_stg_0_28_49, w_stg_0_29_49);
	half_adder ha35( w_stg_1_9_49, w_stg_1_4_50, w_stg_0_30_49, w_stg_0_31_49);
	half_adder ha36( w_stg_1_5_50, w_stg_1_0_51, w_stg_0_19_50, w_stg_0_20_50);
	full_adder_md fa283( w_stg_1_6_50, w_stg_1_1_51, w_stg_0_21_50, w_stg_0_22_50, w_stg_0_23_50);
	full_adder_md fa284( w_stg_1_7_50, w_stg_1_2_51, w_stg_0_24_50, w_stg_0_25_50, w_stg_0_26_50);
	full_adder_md fa285( w_stg_1_8_50, w_stg_1_3_51, w_stg_0_27_50, w_stg_0_28_50, w_stg_0_29_50);
	half_adder ha37( w_stg_1_9_50, w_stg_1_4_51, w_stg_0_30_50, w_stg_0_31_50);
	assign w_stg_1_5_51 = w_stg_0_20_51;
	full_adder_md fa286( w_stg_1_6_51, w_stg_1_0_52, w_stg_0_21_51, w_stg_0_22_51, w_stg_0_23_51);
	full_adder_md fa287( w_stg_1_7_51, w_stg_1_1_52, w_stg_0_24_51, w_stg_0_25_51, w_stg_0_26_51);
	full_adder_md fa288( w_stg_1_8_51, w_stg_1_2_52, w_stg_0_27_51, w_stg_0_28_51, w_stg_0_29_51);
	half_adder ha38( w_stg_1_9_51, w_stg_1_3_52, w_stg_0_30_51, w_stg_0_31_51);
	full_adder_md fa289( w_stg_1_4_52, w_stg_1_0_53, w_stg_0_21_52, w_stg_0_22_52, w_stg_0_23_52);
	full_adder_md fa290( w_stg_1_5_52, w_stg_1_1_53, w_stg_0_24_52, w_stg_0_25_52, w_stg_0_26_52);
	full_adder_md fa291( w_stg_1_6_52, w_stg_1_2_53, w_stg_0_27_52, w_stg_0_28_52, w_stg_0_29_52);
	half_adder ha39( w_stg_1_7_52, w_stg_1_3_53, w_stg_0_30_52, w_stg_0_31_52);
	half_adder ha40( w_stg_1_4_53, w_stg_1_0_54, w_stg_0_22_53, w_stg_0_23_53);
	full_adder_md fa292( w_stg_1_5_53, w_stg_1_1_54, w_stg_0_24_53, w_stg_0_25_53, w_stg_0_26_53);
	full_adder_md fa293( w_stg_1_6_53, w_stg_1_2_54, w_stg_0_27_53, w_stg_0_28_53, w_stg_0_29_53);
	half_adder ha41( w_stg_1_7_53, w_stg_1_3_54, w_stg_0_30_53, w_stg_0_31_53);
	assign w_stg_1_4_54 = w_stg_0_23_54;
	full_adder_md fa294( w_stg_1_5_54, w_stg_1_0_55, w_stg_0_24_54, w_stg_0_25_54, w_stg_0_26_54);
	full_adder_md fa295( w_stg_1_6_54, w_stg_1_1_55, w_stg_0_27_54, w_stg_0_28_54, w_stg_0_29_54);
	half_adder ha42( w_stg_1_7_54, w_stg_1_2_55, w_stg_0_30_54, w_stg_0_31_54);
	full_adder_md fa296( w_stg_1_3_55, w_stg_1_0_56, w_stg_0_24_55, w_stg_0_25_55, w_stg_0_26_55);
	full_adder_md fa297( w_stg_1_4_55, w_stg_1_1_56, w_stg_0_27_55, w_stg_0_28_55, w_stg_0_29_55);
	half_adder ha43( w_stg_1_5_55, w_stg_1_2_56, w_stg_0_30_55, w_stg_0_31_55);
	half_adder ha44( w_stg_1_3_56, w_stg_1_0_57, w_stg_0_25_56, w_stg_0_26_56);
	full_adder_md fa298( w_stg_1_4_56, w_stg_1_1_57, w_stg_0_27_56, w_stg_0_28_56, w_stg_0_29_56);
	half_adder ha45( w_stg_1_5_56, w_stg_1_2_57, w_stg_0_30_56, w_stg_0_31_56);
	assign w_stg_1_3_57 = w_stg_0_26_57;
	full_adder_md fa299( w_stg_1_4_57, w_stg_1_0_58, w_stg_0_27_57, w_stg_0_28_57, w_stg_0_29_57);
	half_adder ha46( w_stg_1_5_57, w_stg_1_1_58, w_stg_0_30_57, w_stg_0_31_57);
	full_adder_md fa300( w_stg_1_2_58, w_stg_1_0_59, w_stg_0_27_58, w_stg_0_28_58, w_stg_0_29_58);
	half_adder ha47( w_stg_1_3_58, w_stg_1_1_59, w_stg_0_30_58, w_stg_0_31_58);
	half_adder ha48( w_stg_1_2_59, w_stg_1_0_60, w_stg_0_28_59, w_stg_0_29_59);
	half_adder ha49( w_stg_1_3_59, w_stg_1_1_60, w_stg_0_30_59, w_stg_0_31_59);
	assign w_stg_1_2_60 = w_stg_0_29_60;
	half_adder ha50( w_stg_1_3_60, w_stg_1_0_61, w_stg_0_30_60, w_stg_0_31_60);
	half_adder ha51( w_stg_1_1_61, w_stg_1_0_62, w_stg_0_30_61, w_stg_0_31_61);
	assign w_stg_1_1_62 = w_stg_0_31_62;
	assign w_stg_2_0_0 = w_stg_1_0_0;
	assign w_stg_2_0_1 = w_stg_1_0_1;
	half_adder ha52( w_stg_2_0_2, w_stg_2_0_3, w_stg_1_0_2, w_stg_1_1_2);
	full_adder_md fa301( w_stg_2_1_3, w_stg_2_0_4, w_stg_1_0_3, w_stg_1_1_3, w_stg_1_2_3);
	full_adder_md fa302( w_stg_2_1_4, w_stg_2_0_5, w_stg_1_0_4, w_stg_1_1_4, w_stg_1_2_4);
	full_adder_md fa303( w_stg_2_1_5, w_stg_2_0_6, w_stg_1_0_5, w_stg_1_1_5, w_stg_1_2_5);
	assign w_stg_2_2_5 = w_stg_1_3_5;
	full_adder_md fa304( w_stg_2_1_6, w_stg_2_0_7, w_stg_1_0_6, w_stg_1_1_6, w_stg_1_2_6);
	half_adder ha53( w_stg_2_2_6, w_stg_2_1_7, w_stg_1_3_6, w_stg_1_4_6);
	full_adder_md fa305( w_stg_2_2_7, w_stg_2_0_8, w_stg_1_0_7, w_stg_1_1_7, w_stg_1_2_7);
	half_adder ha54( w_stg_2_3_7, w_stg_2_1_8, w_stg_1_3_7, w_stg_1_4_7);
	full_adder_md fa306( w_stg_2_2_8, w_stg_2_0_9, w_stg_1_0_8, w_stg_1_1_8, w_stg_1_2_8);
	full_adder_md fa307( w_stg_2_3_8, w_stg_2_1_9, w_stg_1_3_8, w_stg_1_4_8, w_stg_1_5_8);
	full_adder_md fa308( w_stg_2_2_9, w_stg_2_0_10, w_stg_1_0_9, w_stg_1_1_9, w_stg_1_2_9);
	full_adder_md fa309( w_stg_2_3_9, w_stg_2_1_10, w_stg_1_3_9, w_stg_1_4_9, w_stg_1_5_9);
	assign w_stg_2_4_9 = w_stg_1_6_9;
	full_adder_md fa310( w_stg_2_2_10, w_stg_2_0_11, w_stg_1_0_10, w_stg_1_1_10, w_stg_1_2_10);
	full_adder_md fa311( w_stg_2_3_10, w_stg_2_1_11, w_stg_1_3_10, w_stg_1_4_10, w_stg_1_5_10);
	assign w_stg_2_4_10 = w_stg_1_6_10;
	full_adder_md fa312( w_stg_2_2_11, w_stg_2_0_12, w_stg_1_0_11, w_stg_1_1_11, w_stg_1_2_11);
	full_adder_md fa313( w_stg_2_3_11, w_stg_2_1_12, w_stg_1_3_11, w_stg_1_4_11, w_stg_1_5_11);
	half_adder ha55( w_stg_2_4_11, w_stg_2_2_12, w_stg_1_6_11, w_stg_1_7_11);
	full_adder_md fa314( w_stg_2_3_12, w_stg_2_0_13, w_stg_1_0_12, w_stg_1_1_12, w_stg_1_2_12);
	full_adder_md fa315( w_stg_2_4_12, w_stg_2_1_13, w_stg_1_3_12, w_stg_1_4_12, w_stg_1_5_12);
	full_adder_md fa316( w_stg_2_5_12, w_stg_2_2_13, w_stg_1_6_12, w_stg_1_7_12, w_stg_1_8_12);
	full_adder_md fa317( w_stg_2_3_13, w_stg_2_0_14, w_stg_1_0_13, w_stg_1_1_13, w_stg_1_2_13);
	full_adder_md fa318( w_stg_2_4_13, w_stg_2_1_14, w_stg_1_3_13, w_stg_1_4_13, w_stg_1_5_13);
	full_adder_md fa319( w_stg_2_5_13, w_stg_2_2_14, w_stg_1_6_13, w_stg_1_7_13, w_stg_1_8_13);
	full_adder_md fa320( w_stg_2_3_14, w_stg_2_0_15, w_stg_1_0_14, w_stg_1_1_14, w_stg_1_2_14);
	full_adder_md fa321( w_stg_2_4_14, w_stg_2_1_15, w_stg_1_3_14, w_stg_1_4_14, w_stg_1_5_14);
	full_adder_md fa322( w_stg_2_5_14, w_stg_2_2_15, w_stg_1_6_14, w_stg_1_7_14, w_stg_1_8_14);
	assign w_stg_2_6_14 = w_stg_1_9_14;
	full_adder_md fa323( w_stg_2_3_15, w_stg_2_0_16, w_stg_1_0_15, w_stg_1_1_15, w_stg_1_2_15);
	full_adder_md fa324( w_stg_2_4_15, w_stg_2_1_16, w_stg_1_3_15, w_stg_1_4_15, w_stg_1_5_15);
	full_adder_md fa325( w_stg_2_5_15, w_stg_2_2_16, w_stg_1_6_15, w_stg_1_7_15, w_stg_1_8_15);
	half_adder ha56( w_stg_2_6_15, w_stg_2_3_16, w_stg_1_9_15, w_stg_1_10_15);
	full_adder_md fa326( w_stg_2_4_16, w_stg_2_0_17, w_stg_1_0_16, w_stg_1_1_16, w_stg_1_2_16);
	full_adder_md fa327( w_stg_2_5_16, w_stg_2_1_17, w_stg_1_3_16, w_stg_1_4_16, w_stg_1_5_16);
	full_adder_md fa328( w_stg_2_6_16, w_stg_2_2_17, w_stg_1_6_16, w_stg_1_7_16, w_stg_1_8_16);
	half_adder ha57( w_stg_2_7_16, w_stg_2_3_17, w_stg_1_9_16, w_stg_1_10_16);
	full_adder_md fa329( w_stg_2_4_17, w_stg_2_0_18, w_stg_1_0_17, w_stg_1_1_17, w_stg_1_2_17);
	full_adder_md fa330( w_stg_2_5_17, w_stg_2_1_18, w_stg_1_3_17, w_stg_1_4_17, w_stg_1_5_17);
	full_adder_md fa331( w_stg_2_6_17, w_stg_2_2_18, w_stg_1_6_17, w_stg_1_7_17, w_stg_1_8_17);
	full_adder_md fa332( w_stg_2_7_17, w_stg_2_3_18, w_stg_1_9_17, w_stg_1_10_17, w_stg_1_11_17);
	full_adder_md fa333( w_stg_2_4_18, w_stg_2_0_19, w_stg_1_0_18, w_stg_1_1_18, w_stg_1_2_18);
	full_adder_md fa334( w_stg_2_5_18, w_stg_2_1_19, w_stg_1_3_18, w_stg_1_4_18, w_stg_1_5_18);
	full_adder_md fa335( w_stg_2_6_18, w_stg_2_2_19, w_stg_1_6_18, w_stg_1_7_18, w_stg_1_8_18);
	full_adder_md fa336( w_stg_2_7_18, w_stg_2_3_19, w_stg_1_9_18, w_stg_1_10_18, w_stg_1_11_18);
	assign w_stg_2_8_18 = w_stg_1_12_18;
	full_adder_md fa337( w_stg_2_4_19, w_stg_2_0_20, w_stg_1_0_19, w_stg_1_1_19, w_stg_1_2_19);
	full_adder_md fa338( w_stg_2_5_19, w_stg_2_1_20, w_stg_1_3_19, w_stg_1_4_19, w_stg_1_5_19);
	full_adder_md fa339( w_stg_2_6_19, w_stg_2_2_20, w_stg_1_6_19, w_stg_1_7_19, w_stg_1_8_19);
	full_adder_md fa340( w_stg_2_7_19, w_stg_2_3_20, w_stg_1_9_19, w_stg_1_10_19, w_stg_1_11_19);
	assign w_stg_2_8_19 = w_stg_1_12_19;
	full_adder_md fa341( w_stg_2_4_20, w_stg_2_0_21, w_stg_1_0_20, w_stg_1_1_20, w_stg_1_2_20);
	full_adder_md fa342( w_stg_2_5_20, w_stg_2_1_21, w_stg_1_3_20, w_stg_1_4_20, w_stg_1_5_20);
	full_adder_md fa343( w_stg_2_6_20, w_stg_2_2_21, w_stg_1_6_20, w_stg_1_7_20, w_stg_1_8_20);
	full_adder_md fa344( w_stg_2_7_20, w_stg_2_3_21, w_stg_1_9_20, w_stg_1_10_20, w_stg_1_11_20);
	half_adder ha58( w_stg_2_8_20, w_stg_2_4_21, w_stg_1_12_20, w_stg_1_13_20);
	full_adder_md fa345( w_stg_2_5_21, w_stg_2_0_22, w_stg_1_0_21, w_stg_1_1_21, w_stg_1_2_21);
	full_adder_md fa346( w_stg_2_6_21, w_stg_2_1_22, w_stg_1_3_21, w_stg_1_4_21, w_stg_1_5_21);
	full_adder_md fa347( w_stg_2_7_21, w_stg_2_2_22, w_stg_1_6_21, w_stg_1_7_21, w_stg_1_8_21);
	full_adder_md fa348( w_stg_2_8_21, w_stg_2_3_22, w_stg_1_9_21, w_stg_1_10_21, w_stg_1_11_21);
	full_adder_md fa349( w_stg_2_9_21, w_stg_2_4_22, w_stg_1_12_21, w_stg_1_13_21, w_stg_1_14_21);
	full_adder_md fa350( w_stg_2_5_22, w_stg_2_0_23, w_stg_1_0_22, w_stg_1_1_22, w_stg_1_2_22);
	full_adder_md fa351( w_stg_2_6_22, w_stg_2_1_23, w_stg_1_3_22, w_stg_1_4_22, w_stg_1_5_22);
	full_adder_md fa352( w_stg_2_7_22, w_stg_2_2_23, w_stg_1_6_22, w_stg_1_7_22, w_stg_1_8_22);
	full_adder_md fa353( w_stg_2_8_22, w_stg_2_3_23, w_stg_1_9_22, w_stg_1_10_22, w_stg_1_11_22);
	full_adder_md fa354( w_stg_2_9_22, w_stg_2_4_23, w_stg_1_12_22, w_stg_1_13_22, w_stg_1_14_22);
	full_adder_md fa355( w_stg_2_5_23, w_stg_2_0_24, w_stg_1_0_23, w_stg_1_1_23, w_stg_1_2_23);
	full_adder_md fa356( w_stg_2_6_23, w_stg_2_1_24, w_stg_1_3_23, w_stg_1_4_23, w_stg_1_5_23);
	full_adder_md fa357( w_stg_2_7_23, w_stg_2_2_24, w_stg_1_6_23, w_stg_1_7_23, w_stg_1_8_23);
	full_adder_md fa358( w_stg_2_8_23, w_stg_2_3_24, w_stg_1_9_23, w_stg_1_10_23, w_stg_1_11_23);
	full_adder_md fa359( w_stg_2_9_23, w_stg_2_4_24, w_stg_1_12_23, w_stg_1_13_23, w_stg_1_14_23);
	assign w_stg_2_10_23 = w_stg_1_15_23;
	full_adder_md fa360( w_stg_2_5_24, w_stg_2_0_25, w_stg_1_0_24, w_stg_1_1_24, w_stg_1_2_24);
	full_adder_md fa361( w_stg_2_6_24, w_stg_2_1_25, w_stg_1_3_24, w_stg_1_4_24, w_stg_1_5_24);
	full_adder_md fa362( w_stg_2_7_24, w_stg_2_2_25, w_stg_1_6_24, w_stg_1_7_24, w_stg_1_8_24);
	full_adder_md fa363( w_stg_2_8_24, w_stg_2_3_25, w_stg_1_9_24, w_stg_1_10_24, w_stg_1_11_24);
	full_adder_md fa364( w_stg_2_9_24, w_stg_2_4_25, w_stg_1_12_24, w_stg_1_13_24, w_stg_1_14_24);
	half_adder ha59( w_stg_2_10_24, w_stg_2_5_25, w_stg_1_15_24, w_stg_1_16_24);
	full_adder_md fa365( w_stg_2_6_25, w_stg_2_0_26, w_stg_1_0_25, w_stg_1_1_25, w_stg_1_2_25);
	full_adder_md fa366( w_stg_2_7_25, w_stg_2_1_26, w_stg_1_3_25, w_stg_1_4_25, w_stg_1_5_25);
	full_adder_md fa367( w_stg_2_8_25, w_stg_2_2_26, w_stg_1_6_25, w_stg_1_7_25, w_stg_1_8_25);
	full_adder_md fa368( w_stg_2_9_25, w_stg_2_3_26, w_stg_1_9_25, w_stg_1_10_25, w_stg_1_11_25);
	full_adder_md fa369( w_stg_2_10_25, w_stg_2_4_26, w_stg_1_12_25, w_stg_1_13_25, w_stg_1_14_25);
	half_adder ha60( w_stg_2_11_25, w_stg_2_5_26, w_stg_1_15_25, w_stg_1_16_25);
	full_adder_md fa370( w_stg_2_6_26, w_stg_2_0_27, w_stg_1_0_26, w_stg_1_1_26, w_stg_1_2_26);
	full_adder_md fa371( w_stg_2_7_26, w_stg_2_1_27, w_stg_1_3_26, w_stg_1_4_26, w_stg_1_5_26);
	full_adder_md fa372( w_stg_2_8_26, w_stg_2_2_27, w_stg_1_6_26, w_stg_1_7_26, w_stg_1_8_26);
	full_adder_md fa373( w_stg_2_9_26, w_stg_2_3_27, w_stg_1_9_26, w_stg_1_10_26, w_stg_1_11_26);
	full_adder_md fa374( w_stg_2_10_26, w_stg_2_4_27, w_stg_1_12_26, w_stg_1_13_26, w_stg_1_14_26);
	full_adder_md fa375( w_stg_2_11_26, w_stg_2_5_27, w_stg_1_15_26, w_stg_1_16_26, w_stg_1_17_26);
	full_adder_md fa376( w_stg_2_6_27, w_stg_2_0_28, w_stg_1_0_27, w_stg_1_1_27, w_stg_1_2_27);
	full_adder_md fa377( w_stg_2_7_27, w_stg_2_1_28, w_stg_1_3_27, w_stg_1_4_27, w_stg_1_5_27);
	full_adder_md fa378( w_stg_2_8_27, w_stg_2_2_28, w_stg_1_6_27, w_stg_1_7_27, w_stg_1_8_27);
	full_adder_md fa379( w_stg_2_9_27, w_stg_2_3_28, w_stg_1_9_27, w_stg_1_10_27, w_stg_1_11_27);
	full_adder_md fa380( w_stg_2_10_27, w_stg_2_4_28, w_stg_1_12_27, w_stg_1_13_27, w_stg_1_14_27);
	full_adder_md fa381( w_stg_2_11_27, w_stg_2_5_28, w_stg_1_15_27, w_stg_1_16_27, w_stg_1_17_27);
	assign w_stg_2_12_27 = w_stg_1_18_27;
	full_adder_md fa382( w_stg_2_6_28, w_stg_2_0_29, w_stg_1_0_28, w_stg_1_1_28, w_stg_1_2_28);
	full_adder_md fa383( w_stg_2_7_28, w_stg_2_1_29, w_stg_1_3_28, w_stg_1_4_28, w_stg_1_5_28);
	full_adder_md fa384( w_stg_2_8_28, w_stg_2_2_29, w_stg_1_6_28, w_stg_1_7_28, w_stg_1_8_28);
	full_adder_md fa385( w_stg_2_9_28, w_stg_2_3_29, w_stg_1_9_28, w_stg_1_10_28, w_stg_1_11_28);
	full_adder_md fa386( w_stg_2_10_28, w_stg_2_4_29, w_stg_1_12_28, w_stg_1_13_28, w_stg_1_14_28);
	full_adder_md fa387( w_stg_2_11_28, w_stg_2_5_29, w_stg_1_15_28, w_stg_1_16_28, w_stg_1_17_28);
	assign w_stg_2_12_28 = w_stg_1_18_28;
	full_adder_md fa388( w_stg_2_6_29, w_stg_2_0_30, w_stg_1_0_29, w_stg_1_1_29, w_stg_1_2_29);
	full_adder_md fa389( w_stg_2_7_29, w_stg_2_1_30, w_stg_1_3_29, w_stg_1_4_29, w_stg_1_5_29);
	full_adder_md fa390( w_stg_2_8_29, w_stg_2_2_30, w_stg_1_6_29, w_stg_1_7_29, w_stg_1_8_29);
	full_adder_md fa391( w_stg_2_9_29, w_stg_2_3_30, w_stg_1_9_29, w_stg_1_10_29, w_stg_1_11_29);
	full_adder_md fa392( w_stg_2_10_29, w_stg_2_4_30, w_stg_1_12_29, w_stg_1_13_29, w_stg_1_14_29);
	full_adder_md fa393( w_stg_2_11_29, w_stg_2_5_30, w_stg_1_15_29, w_stg_1_16_29, w_stg_1_17_29);
	half_adder ha61( w_stg_2_12_29, w_stg_2_6_30, w_stg_1_18_29, w_stg_1_19_29);
	full_adder_md fa394( w_stg_2_7_30, w_stg_2_0_31, w_stg_1_0_30, w_stg_1_1_30, w_stg_1_2_30);
	full_adder_md fa395( w_stg_2_8_30, w_stg_2_1_31, w_stg_1_3_30, w_stg_1_4_30, w_stg_1_5_30);
	full_adder_md fa396( w_stg_2_9_30, w_stg_2_2_31, w_stg_1_6_30, w_stg_1_7_30, w_stg_1_8_30);
	full_adder_md fa397( w_stg_2_10_30, w_stg_2_3_31, w_stg_1_9_30, w_stg_1_10_30, w_stg_1_11_30);
	full_adder_md fa398( w_stg_2_11_30, w_stg_2_4_31, w_stg_1_12_30, w_stg_1_13_30, w_stg_1_14_30);
	full_adder_md fa399( w_stg_2_12_30, w_stg_2_5_31, w_stg_1_15_30, w_stg_1_16_30, w_stg_1_17_30);
	full_adder_md fa400( w_stg_2_13_30, w_stg_2_6_31, w_stg_1_18_30, w_stg_1_19_30, w_stg_1_20_30);
	full_adder_md fa401( w_stg_2_7_31, w_stg_2_0_32, w_stg_1_0_31, w_stg_1_1_31, w_stg_1_2_31);
	full_adder_md fa402( w_stg_2_8_31, w_stg_2_1_32, w_stg_1_3_31, w_stg_1_4_31, w_stg_1_5_31);
	full_adder_md fa403( w_stg_2_9_31, w_stg_2_2_32, w_stg_1_6_31, w_stg_1_7_31, w_stg_1_8_31);
	full_adder_md fa404( w_stg_2_10_31, w_stg_2_3_32, w_stg_1_9_31, w_stg_1_10_31, w_stg_1_11_31);
	full_adder_md fa405( w_stg_2_11_31, w_stg_2_4_32, w_stg_1_12_31, w_stg_1_13_31, w_stg_1_14_31);
	full_adder_md fa406( w_stg_2_12_31, w_stg_2_5_32, w_stg_1_15_31, w_stg_1_16_31, w_stg_1_17_31);
	full_adder_md fa407( w_stg_2_13_31, w_stg_2_6_32, w_stg_1_18_31, w_stg_1_19_31, w_stg_1_20_31);
	full_adder_md fa408( w_stg_2_7_32, w_stg_2_0_33, w_stg_1_0_32, w_stg_1_1_32, w_stg_1_2_32);
	full_adder_md fa409( w_stg_2_8_32, w_stg_2_1_33, w_stg_1_3_32, w_stg_1_4_32, w_stg_1_5_32);
	full_adder_md fa410( w_stg_2_9_32, w_stg_2_2_33, w_stg_1_6_32, w_stg_1_7_32, w_stg_1_8_32);
	full_adder_md fa411( w_stg_2_10_32, w_stg_2_3_33, w_stg_1_9_32, w_stg_1_10_32, w_stg_1_11_32);
	full_adder_md fa412( w_stg_2_11_32, w_stg_2_4_33, w_stg_1_12_32, w_stg_1_13_32, w_stg_1_14_32);
	full_adder_md fa413( w_stg_2_12_32, w_stg_2_5_33, w_stg_1_15_32, w_stg_1_16_32, w_stg_1_17_32);
	full_adder_md fa414( w_stg_2_13_32, w_stg_2_6_33, w_stg_1_18_32, w_stg_1_19_32, w_stg_1_20_32);
	assign w_stg_2_14_32 = w_stg_1_21_32;
	full_adder_md fa415( w_stg_2_7_33, w_stg_2_0_34, w_stg_1_0_33, w_stg_1_1_33, w_stg_1_2_33);
	full_adder_md fa416( w_stg_2_8_33, w_stg_2_1_34, w_stg_1_3_33, w_stg_1_4_33, w_stg_1_5_33);
	full_adder_md fa417( w_stg_2_9_33, w_stg_2_2_34, w_stg_1_6_33, w_stg_1_7_33, w_stg_1_8_33);
	full_adder_md fa418( w_stg_2_10_33, w_stg_2_3_34, w_stg_1_9_33, w_stg_1_10_33, w_stg_1_11_33);
	full_adder_md fa419( w_stg_2_11_33, w_stg_2_4_34, w_stg_1_12_33, w_stg_1_13_33, w_stg_1_14_33);
	full_adder_md fa420( w_stg_2_12_33, w_stg_2_5_34, w_stg_1_15_33, w_stg_1_16_33, w_stg_1_17_33);
	full_adder_md fa421( w_stg_2_13_33, w_stg_2_6_34, w_stg_1_18_33, w_stg_1_19_33, w_stg_1_20_33);
	assign w_stg_2_14_33 = w_stg_1_21_33;
	full_adder_md fa422( w_stg_2_7_34, w_stg_2_0_35, w_stg_1_0_34, w_stg_1_1_34, w_stg_1_2_34);
	full_adder_md fa423( w_stg_2_8_34, w_stg_2_1_35, w_stg_1_3_34, w_stg_1_4_34, w_stg_1_5_34);
	full_adder_md fa424( w_stg_2_9_34, w_stg_2_2_35, w_stg_1_6_34, w_stg_1_7_34, w_stg_1_8_34);
	full_adder_md fa425( w_stg_2_10_34, w_stg_2_3_35, w_stg_1_9_34, w_stg_1_10_34, w_stg_1_11_34);
	full_adder_md fa426( w_stg_2_11_34, w_stg_2_4_35, w_stg_1_12_34, w_stg_1_13_34, w_stg_1_14_34);
	full_adder_md fa427( w_stg_2_12_34, w_stg_2_5_35, w_stg_1_15_34, w_stg_1_16_34, w_stg_1_17_34);
	half_adder ha62( w_stg_2_13_34, w_stg_2_6_35, w_stg_1_18_34, w_stg_1_19_34);
	full_adder_md fa428( w_stg_2_7_35, w_stg_2_0_36, w_stg_1_0_35, w_stg_1_1_35, w_stg_1_2_35);
	full_adder_md fa429( w_stg_2_8_35, w_stg_2_1_36, w_stg_1_3_35, w_stg_1_4_35, w_stg_1_5_35);
	full_adder_md fa430( w_stg_2_9_35, w_stg_2_2_36, w_stg_1_6_35, w_stg_1_7_35, w_stg_1_8_35);
	full_adder_md fa431( w_stg_2_10_35, w_stg_2_3_36, w_stg_1_9_35, w_stg_1_10_35, w_stg_1_11_35);
	full_adder_md fa432( w_stg_2_11_35, w_stg_2_4_36, w_stg_1_12_35, w_stg_1_13_35, w_stg_1_14_35);
	full_adder_md fa433( w_stg_2_12_35, w_stg_2_5_36, w_stg_1_15_35, w_stg_1_16_35, w_stg_1_17_35);
	half_adder ha63( w_stg_2_13_35, w_stg_2_6_36, w_stg_1_18_35, w_stg_1_19_35);
	full_adder_md fa434( w_stg_2_7_36, w_stg_2_0_37, w_stg_1_0_36, w_stg_1_1_36, w_stg_1_2_36);
	full_adder_md fa435( w_stg_2_8_36, w_stg_2_1_37, w_stg_1_3_36, w_stg_1_4_36, w_stg_1_5_36);
	full_adder_md fa436( w_stg_2_9_36, w_stg_2_2_37, w_stg_1_6_36, w_stg_1_7_36, w_stg_1_8_36);
	full_adder_md fa437( w_stg_2_10_36, w_stg_2_3_37, w_stg_1_9_36, w_stg_1_10_36, w_stg_1_11_36);
	full_adder_md fa438( w_stg_2_11_36, w_stg_2_4_37, w_stg_1_12_36, w_stg_1_13_36, w_stg_1_14_36);
	full_adder_md fa439( w_stg_2_12_36, w_stg_2_5_37, w_stg_1_15_36, w_stg_1_16_36, w_stg_1_17_36);
	half_adder ha64( w_stg_2_13_36, w_stg_2_6_37, w_stg_1_18_36, w_stg_1_19_36);
	full_adder_md fa440( w_stg_2_7_37, w_stg_2_0_38, w_stg_1_0_37, w_stg_1_1_37, w_stg_1_2_37);
	full_adder_md fa441( w_stg_2_8_37, w_stg_2_1_38, w_stg_1_3_37, w_stg_1_4_37, w_stg_1_5_37);
	full_adder_md fa442( w_stg_2_9_37, w_stg_2_2_38, w_stg_1_6_37, w_stg_1_7_37, w_stg_1_8_37);
	full_adder_md fa443( w_stg_2_10_37, w_stg_2_3_38, w_stg_1_9_37, w_stg_1_10_37, w_stg_1_11_37);
	full_adder_md fa444( w_stg_2_11_37, w_stg_2_4_38, w_stg_1_12_37, w_stg_1_13_37, w_stg_1_14_37);
	full_adder_md fa445( w_stg_2_12_37, w_stg_2_5_38, w_stg_1_15_37, w_stg_1_16_37, w_stg_1_17_37);
	full_adder_md fa446( w_stg_2_6_38, w_stg_2_0_39, w_stg_1_0_38, w_stg_1_1_38, w_stg_1_2_38);
	full_adder_md fa447( w_stg_2_7_38, w_stg_2_1_39, w_stg_1_3_38, w_stg_1_4_38, w_stg_1_5_38);
	full_adder_md fa448( w_stg_2_8_38, w_stg_2_2_39, w_stg_1_6_38, w_stg_1_7_38, w_stg_1_8_38);
	full_adder_md fa449( w_stg_2_9_38, w_stg_2_3_39, w_stg_1_9_38, w_stg_1_10_38, w_stg_1_11_38);
	full_adder_md fa450( w_stg_2_10_38, w_stg_2_4_39, w_stg_1_12_38, w_stg_1_13_38, w_stg_1_14_38);
	full_adder_md fa451( w_stg_2_11_38, w_stg_2_5_39, w_stg_1_15_38, w_stg_1_16_38, w_stg_1_17_38);
	full_adder_md fa452( w_stg_2_6_39, w_stg_2_0_40, w_stg_1_0_39, w_stg_1_1_39, w_stg_1_2_39);
	full_adder_md fa453( w_stg_2_7_39, w_stg_2_1_40, w_stg_1_3_39, w_stg_1_4_39, w_stg_1_5_39);
	full_adder_md fa454( w_stg_2_8_39, w_stg_2_2_40, w_stg_1_6_39, w_stg_1_7_39, w_stg_1_8_39);
	full_adder_md fa455( w_stg_2_9_39, w_stg_2_3_40, w_stg_1_9_39, w_stg_1_10_39, w_stg_1_11_39);
	full_adder_md fa456( w_stg_2_10_39, w_stg_2_4_40, w_stg_1_12_39, w_stg_1_13_39, w_stg_1_14_39);
	full_adder_md fa457( w_stg_2_11_39, w_stg_2_5_40, w_stg_1_15_39, w_stg_1_16_39, w_stg_1_17_39);
	full_adder_md fa458( w_stg_2_6_40, w_stg_2_0_41, w_stg_1_0_40, w_stg_1_1_40, w_stg_1_2_40);
	full_adder_md fa459( w_stg_2_7_40, w_stg_2_1_41, w_stg_1_3_40, w_stg_1_4_40, w_stg_1_5_40);
	full_adder_md fa460( w_stg_2_8_40, w_stg_2_2_41, w_stg_1_6_40, w_stg_1_7_40, w_stg_1_8_40);
	full_adder_md fa461( w_stg_2_9_40, w_stg_2_3_41, w_stg_1_9_40, w_stg_1_10_40, w_stg_1_11_40);
	full_adder_md fa462( w_stg_2_10_40, w_stg_2_4_41, w_stg_1_12_40, w_stg_1_13_40, w_stg_1_14_40);
	assign w_stg_2_11_40 = w_stg_1_15_40;
	full_adder_md fa463( w_stg_2_5_41, w_stg_2_0_42, w_stg_1_0_41, w_stg_1_1_41, w_stg_1_2_41);
	full_adder_md fa464( w_stg_2_6_41, w_stg_2_1_42, w_stg_1_3_41, w_stg_1_4_41, w_stg_1_5_41);
	full_adder_md fa465( w_stg_2_7_41, w_stg_2_2_42, w_stg_1_6_41, w_stg_1_7_41, w_stg_1_8_41);
	full_adder_md fa466( w_stg_2_8_41, w_stg_2_3_42, w_stg_1_9_41, w_stg_1_10_41, w_stg_1_11_41);
	full_adder_md fa467( w_stg_2_9_41, w_stg_2_4_42, w_stg_1_12_41, w_stg_1_13_41, w_stg_1_14_41);
	assign w_stg_2_10_41 = w_stg_1_15_41;
	full_adder_md fa468( w_stg_2_5_42, w_stg_2_0_43, w_stg_1_0_42, w_stg_1_1_42, w_stg_1_2_42);
	full_adder_md fa469( w_stg_2_6_42, w_stg_2_1_43, w_stg_1_3_42, w_stg_1_4_42, w_stg_1_5_42);
	full_adder_md fa470( w_stg_2_7_42, w_stg_2_2_43, w_stg_1_6_42, w_stg_1_7_42, w_stg_1_8_42);
	full_adder_md fa471( w_stg_2_8_42, w_stg_2_3_43, w_stg_1_9_42, w_stg_1_10_42, w_stg_1_11_42);
	full_adder_md fa472( w_stg_2_9_42, w_stg_2_4_43, w_stg_1_12_42, w_stg_1_13_42, w_stg_1_14_42);
	assign w_stg_2_10_42 = w_stg_1_15_42;
	full_adder_md fa473( w_stg_2_5_43, w_stg_2_0_44, w_stg_1_0_43, w_stg_1_1_43, w_stg_1_2_43);
	full_adder_md fa474( w_stg_2_6_43, w_stg_2_1_44, w_stg_1_3_43, w_stg_1_4_43, w_stg_1_5_43);
	full_adder_md fa475( w_stg_2_7_43, w_stg_2_2_44, w_stg_1_6_43, w_stg_1_7_43, w_stg_1_8_43);
	full_adder_md fa476( w_stg_2_8_43, w_stg_2_3_44, w_stg_1_9_43, w_stg_1_10_43, w_stg_1_11_43);
	half_adder ha65( w_stg_2_9_43, w_stg_2_4_44, w_stg_1_12_43, w_stg_1_13_43);
	full_adder_md fa477( w_stg_2_5_44, w_stg_2_0_45, w_stg_1_0_44, w_stg_1_1_44, w_stg_1_2_44);
	full_adder_md fa478( w_stg_2_6_44, w_stg_2_1_45, w_stg_1_3_44, w_stg_1_4_44, w_stg_1_5_44);
	full_adder_md fa479( w_stg_2_7_44, w_stg_2_2_45, w_stg_1_6_44, w_stg_1_7_44, w_stg_1_8_44);
	full_adder_md fa480( w_stg_2_8_44, w_stg_2_3_45, w_stg_1_9_44, w_stg_1_10_44, w_stg_1_11_44);
	half_adder ha66( w_stg_2_9_44, w_stg_2_4_45, w_stg_1_12_44, w_stg_1_13_44);
	full_adder_md fa481( w_stg_2_5_45, w_stg_2_0_46, w_stg_1_0_45, w_stg_1_1_45, w_stg_1_2_45);
	full_adder_md fa482( w_stg_2_6_45, w_stg_2_1_46, w_stg_1_3_45, w_stg_1_4_45, w_stg_1_5_45);
	full_adder_md fa483( w_stg_2_7_45, w_stg_2_2_46, w_stg_1_6_45, w_stg_1_7_45, w_stg_1_8_45);
	full_adder_md fa484( w_stg_2_8_45, w_stg_2_3_46, w_stg_1_9_45, w_stg_1_10_45, w_stg_1_11_45);
	half_adder ha67( w_stg_2_9_45, w_stg_2_4_46, w_stg_1_12_45, w_stg_1_13_45);
	full_adder_md fa485( w_stg_2_5_46, w_stg_2_0_47, w_stg_1_0_46, w_stg_1_1_46, w_stg_1_2_46);
	full_adder_md fa486( w_stg_2_6_46, w_stg_2_1_47, w_stg_1_3_46, w_stg_1_4_46, w_stg_1_5_46);
	full_adder_md fa487( w_stg_2_7_46, w_stg_2_2_47, w_stg_1_6_46, w_stg_1_7_46, w_stg_1_8_46);
	full_adder_md fa488( w_stg_2_8_46, w_stg_2_3_47, w_stg_1_9_46, w_stg_1_10_46, w_stg_1_11_46);
	full_adder_md fa489( w_stg_2_4_47, w_stg_2_0_48, w_stg_1_0_47, w_stg_1_1_47, w_stg_1_2_47);
	full_adder_md fa490( w_stg_2_5_47, w_stg_2_1_48, w_stg_1_3_47, w_stg_1_4_47, w_stg_1_5_47);
	full_adder_md fa491( w_stg_2_6_47, w_stg_2_2_48, w_stg_1_6_47, w_stg_1_7_47, w_stg_1_8_47);
	full_adder_md fa492( w_stg_2_7_47, w_stg_2_3_48, w_stg_1_9_47, w_stg_1_10_47, w_stg_1_11_47);
	full_adder_md fa493( w_stg_2_4_48, w_stg_2_0_49, w_stg_1_0_48, w_stg_1_1_48, w_stg_1_2_48);
	full_adder_md fa494( w_stg_2_5_48, w_stg_2_1_49, w_stg_1_3_48, w_stg_1_4_48, w_stg_1_5_48);
	full_adder_md fa495( w_stg_2_6_48, w_stg_2_2_49, w_stg_1_6_48, w_stg_1_7_48, w_stg_1_8_48);
	full_adder_md fa496( w_stg_2_7_48, w_stg_2_3_49, w_stg_1_9_48, w_stg_1_10_48, w_stg_1_11_48);
	full_adder_md fa497( w_stg_2_4_49, w_stg_2_0_50, w_stg_1_0_49, w_stg_1_1_49, w_stg_1_2_49);
	full_adder_md fa498( w_stg_2_5_49, w_stg_2_1_50, w_stg_1_3_49, w_stg_1_4_49, w_stg_1_5_49);
	full_adder_md fa499( w_stg_2_6_49, w_stg_2_2_50, w_stg_1_6_49, w_stg_1_7_49, w_stg_1_8_49);
	assign w_stg_2_7_49 = w_stg_1_9_49;
	full_adder_md fa500( w_stg_2_3_50, w_stg_2_0_51, w_stg_1_0_50, w_stg_1_1_50, w_stg_1_2_50);
	full_adder_md fa501( w_stg_2_4_50, w_stg_2_1_51, w_stg_1_3_50, w_stg_1_4_50, w_stg_1_5_50);
	full_adder_md fa502( w_stg_2_5_50, w_stg_2_2_51, w_stg_1_6_50, w_stg_1_7_50, w_stg_1_8_50);
	assign w_stg_2_6_50 = w_stg_1_9_50;
	full_adder_md fa503( w_stg_2_3_51, w_stg_2_0_52, w_stg_1_0_51, w_stg_1_1_51, w_stg_1_2_51);
	full_adder_md fa504( w_stg_2_4_51, w_stg_2_1_52, w_stg_1_3_51, w_stg_1_4_51, w_stg_1_5_51);
	full_adder_md fa505( w_stg_2_5_51, w_stg_2_2_52, w_stg_1_6_51, w_stg_1_7_51, w_stg_1_8_51);
	assign w_stg_2_6_51 = w_stg_1_9_51;
	full_adder_md fa506( w_stg_2_3_52, w_stg_2_0_53, w_stg_1_0_52, w_stg_1_1_52, w_stg_1_2_52);
	full_adder_md fa507( w_stg_2_4_52, w_stg_2_1_53, w_stg_1_3_52, w_stg_1_4_52, w_stg_1_5_52);
	half_adder ha68( w_stg_2_5_52, w_stg_2_2_53, w_stg_1_6_52, w_stg_1_7_52);
	full_adder_md fa508( w_stg_2_3_53, w_stg_2_0_54, w_stg_1_0_53, w_stg_1_1_53, w_stg_1_2_53);
	full_adder_md fa509( w_stg_2_4_53, w_stg_2_1_54, w_stg_1_3_53, w_stg_1_4_53, w_stg_1_5_53);
	half_adder ha69( w_stg_2_5_53, w_stg_2_2_54, w_stg_1_6_53, w_stg_1_7_53);
	full_adder_md fa510( w_stg_2_3_54, w_stg_2_0_55, w_stg_1_0_54, w_stg_1_1_54, w_stg_1_2_54);
	full_adder_md fa511( w_stg_2_4_54, w_stg_2_1_55, w_stg_1_3_54, w_stg_1_4_54, w_stg_1_5_54);
	half_adder ha70( w_stg_2_5_54, w_stg_2_2_55, w_stg_1_6_54, w_stg_1_7_54);
	full_adder_md fa512( w_stg_2_3_55, w_stg_2_0_56, w_stg_1_0_55, w_stg_1_1_55, w_stg_1_2_55);
	full_adder_md fa513( w_stg_2_4_55, w_stg_2_1_56, w_stg_1_3_55, w_stg_1_4_55, w_stg_1_5_55);
	full_adder_md fa514( w_stg_2_2_56, w_stg_2_0_57, w_stg_1_0_56, w_stg_1_1_56, w_stg_1_2_56);
	full_adder_md fa515( w_stg_2_3_56, w_stg_2_1_57, w_stg_1_3_56, w_stg_1_4_56, w_stg_1_5_56);
	full_adder_md fa516( w_stg_2_2_57, w_stg_2_0_58, w_stg_1_0_57, w_stg_1_1_57, w_stg_1_2_57);
	full_adder_md fa517( w_stg_2_3_57, w_stg_2_1_58, w_stg_1_3_57, w_stg_1_4_57, w_stg_1_5_57);
	full_adder_md fa518( w_stg_2_2_58, w_stg_2_0_59, w_stg_1_0_58, w_stg_1_1_58, w_stg_1_2_58);
	assign w_stg_2_3_58 = w_stg_1_3_58;
	full_adder_md fa519( w_stg_2_1_59, w_stg_2_0_60, w_stg_1_0_59, w_stg_1_1_59, w_stg_1_2_59);
	assign w_stg_2_2_59 = w_stg_1_3_59;
	full_adder_md fa520( w_stg_2_1_60, w_stg_2_0_61, w_stg_1_0_60, w_stg_1_1_60, w_stg_1_2_60);
	assign w_stg_2_2_60 = w_stg_1_3_60;
	half_adder ha71( w_stg_2_1_61, w_stg_2_0_62, w_stg_1_0_61, w_stg_1_1_61);
	half_adder ha72( w_stg_2_1_62, w_stg_2_0_63, w_stg_1_0_62, w_stg_1_1_62);
	assign w_stg_3_0_0 = w_stg_2_0_0;
	assign w_stg_3_0_1 = w_stg_2_0_1;
	assign w_stg_3_0_2 = w_stg_2_0_2;
	half_adder ha73( w_stg_3_0_3, w_stg_3_0_4, w_stg_2_0_3, w_stg_2_1_3);
	half_adder ha74( w_stg_3_1_4, w_stg_3_0_5, w_stg_2_0_4, w_stg_2_1_4);
	full_adder_md fa521( w_stg_3_1_5, w_stg_3_0_6, w_stg_2_0_5, w_stg_2_1_5, w_stg_2_2_5);
	full_adder_md fa522( w_stg_3_1_6, w_stg_3_0_7, w_stg_2_0_6, w_stg_2_1_6, w_stg_2_2_6);
	full_adder_md fa523( w_stg_3_1_7, w_stg_3_0_8, w_stg_2_0_7, w_stg_2_1_7, w_stg_2_2_7);
	assign w_stg_3_2_7 = w_stg_2_3_7;
	full_adder_md fa524( w_stg_3_1_8, w_stg_3_0_9, w_stg_2_0_8, w_stg_2_1_8, w_stg_2_2_8);
	assign w_stg_3_2_8 = w_stg_2_3_8;
	full_adder_md fa525( w_stg_3_1_9, w_stg_3_0_10, w_stg_2_0_9, w_stg_2_1_9, w_stg_2_2_9);
	half_adder ha75( w_stg_3_2_9, w_stg_3_1_10, w_stg_2_3_9, w_stg_2_4_9);
	full_adder_md fa526( w_stg_3_2_10, w_stg_3_0_11, w_stg_2_0_10, w_stg_2_1_10, w_stg_2_2_10);
	half_adder ha76( w_stg_3_3_10, w_stg_3_1_11, w_stg_2_3_10, w_stg_2_4_10);
	full_adder_md fa527( w_stg_3_2_11, w_stg_3_0_12, w_stg_2_0_11, w_stg_2_1_11, w_stg_2_2_11);
	half_adder ha77( w_stg_3_3_11, w_stg_3_1_12, w_stg_2_3_11, w_stg_2_4_11);
	full_adder_md fa528( w_stg_3_2_12, w_stg_3_0_13, w_stg_2_0_12, w_stg_2_1_12, w_stg_2_2_12);
	full_adder_md fa529( w_stg_3_3_12, w_stg_3_1_13, w_stg_2_3_12, w_stg_2_4_12, w_stg_2_5_12);
	full_adder_md fa530( w_stg_3_2_13, w_stg_3_0_14, w_stg_2_0_13, w_stg_2_1_13, w_stg_2_2_13);
	full_adder_md fa531( w_stg_3_3_13, w_stg_3_1_14, w_stg_2_3_13, w_stg_2_4_13, w_stg_2_5_13);
	full_adder_md fa532( w_stg_3_2_14, w_stg_3_0_15, w_stg_2_0_14, w_stg_2_1_14, w_stg_2_2_14);
	full_adder_md fa533( w_stg_3_3_14, w_stg_3_1_15, w_stg_2_3_14, w_stg_2_4_14, w_stg_2_5_14);
	assign w_stg_3_4_14 = w_stg_2_6_14;
	full_adder_md fa534( w_stg_3_2_15, w_stg_3_0_16, w_stg_2_0_15, w_stg_2_1_15, w_stg_2_2_15);
	full_adder_md fa535( w_stg_3_3_15, w_stg_3_1_16, w_stg_2_3_15, w_stg_2_4_15, w_stg_2_5_15);
	assign w_stg_3_4_15 = w_stg_2_6_15;
	full_adder_md fa536( w_stg_3_2_16, w_stg_3_0_17, w_stg_2_0_16, w_stg_2_1_16, w_stg_2_2_16);
	full_adder_md fa537( w_stg_3_3_16, w_stg_3_1_17, w_stg_2_3_16, w_stg_2_4_16, w_stg_2_5_16);
	half_adder ha78( w_stg_3_4_16, w_stg_3_2_17, w_stg_2_6_16, w_stg_2_7_16);
	full_adder_md fa538( w_stg_3_3_17, w_stg_3_0_18, w_stg_2_0_17, w_stg_2_1_17, w_stg_2_2_17);
	full_adder_md fa539( w_stg_3_4_17, w_stg_3_1_18, w_stg_2_3_17, w_stg_2_4_17, w_stg_2_5_17);
	half_adder ha79( w_stg_3_5_17, w_stg_3_2_18, w_stg_2_6_17, w_stg_2_7_17);
	full_adder_md fa540( w_stg_3_3_18, w_stg_3_0_19, w_stg_2_0_18, w_stg_2_1_18, w_stg_2_2_18);
	full_adder_md fa541( w_stg_3_4_18, w_stg_3_1_19, w_stg_2_3_18, w_stg_2_4_18, w_stg_2_5_18);
	full_adder_md fa542( w_stg_3_5_18, w_stg_3_2_19, w_stg_2_6_18, w_stg_2_7_18, w_stg_2_8_18);
	full_adder_md fa543( w_stg_3_3_19, w_stg_3_0_20, w_stg_2_0_19, w_stg_2_1_19, w_stg_2_2_19);
	full_adder_md fa544( w_stg_3_4_19, w_stg_3_1_20, w_stg_2_3_19, w_stg_2_4_19, w_stg_2_5_19);
	full_adder_md fa545( w_stg_3_5_19, w_stg_3_2_20, w_stg_2_6_19, w_stg_2_7_19, w_stg_2_8_19);
	full_adder_md fa546( w_stg_3_3_20, w_stg_3_0_21, w_stg_2_0_20, w_stg_2_1_20, w_stg_2_2_20);
	full_adder_md fa547( w_stg_3_4_20, w_stg_3_1_21, w_stg_2_3_20, w_stg_2_4_20, w_stg_2_5_20);
	full_adder_md fa548( w_stg_3_5_20, w_stg_3_2_21, w_stg_2_6_20, w_stg_2_7_20, w_stg_2_8_20);
	full_adder_md fa549( w_stg_3_3_21, w_stg_3_0_22, w_stg_2_0_21, w_stg_2_1_21, w_stg_2_2_21);
	full_adder_md fa550( w_stg_3_4_21, w_stg_3_1_22, w_stg_2_3_21, w_stg_2_4_21, w_stg_2_5_21);
	full_adder_md fa551( w_stg_3_5_21, w_stg_3_2_22, w_stg_2_6_21, w_stg_2_7_21, w_stg_2_8_21);
	assign w_stg_3_6_21 = w_stg_2_9_21;
	full_adder_md fa552( w_stg_3_3_22, w_stg_3_0_23, w_stg_2_0_22, w_stg_2_1_22, w_stg_2_2_22);
	full_adder_md fa553( w_stg_3_4_22, w_stg_3_1_23, w_stg_2_3_22, w_stg_2_4_22, w_stg_2_5_22);
	full_adder_md fa554( w_stg_3_5_22, w_stg_3_2_23, w_stg_2_6_22, w_stg_2_7_22, w_stg_2_8_22);
	assign w_stg_3_6_22 = w_stg_2_9_22;
	full_adder_md fa555( w_stg_3_3_23, w_stg_3_0_24, w_stg_2_0_23, w_stg_2_1_23, w_stg_2_2_23);
	full_adder_md fa556( w_stg_3_4_23, w_stg_3_1_24, w_stg_2_3_23, w_stg_2_4_23, w_stg_2_5_23);
	full_adder_md fa557( w_stg_3_5_23, w_stg_3_2_24, w_stg_2_6_23, w_stg_2_7_23, w_stg_2_8_23);
	half_adder ha80( w_stg_3_6_23, w_stg_3_3_24, w_stg_2_9_23, w_stg_2_10_23);
	full_adder_md fa558( w_stg_3_4_24, w_stg_3_0_25, w_stg_2_0_24, w_stg_2_1_24, w_stg_2_2_24);
	full_adder_md fa559( w_stg_3_5_24, w_stg_3_1_25, w_stg_2_3_24, w_stg_2_4_24, w_stg_2_5_24);
	full_adder_md fa560( w_stg_3_6_24, w_stg_3_2_25, w_stg_2_6_24, w_stg_2_7_24, w_stg_2_8_24);
	half_adder ha81( w_stg_3_7_24, w_stg_3_3_25, w_stg_2_9_24, w_stg_2_10_24);
	full_adder_md fa561( w_stg_3_4_25, w_stg_3_0_26, w_stg_2_0_25, w_stg_2_1_25, w_stg_2_2_25);
	full_adder_md fa562( w_stg_3_5_25, w_stg_3_1_26, w_stg_2_3_25, w_stg_2_4_25, w_stg_2_5_25);
	full_adder_md fa563( w_stg_3_6_25, w_stg_3_2_26, w_stg_2_6_25, w_stg_2_7_25, w_stg_2_8_25);
	full_adder_md fa564( w_stg_3_7_25, w_stg_3_3_26, w_stg_2_9_25, w_stg_2_10_25, w_stg_2_11_25);
	full_adder_md fa565( w_stg_3_4_26, w_stg_3_0_27, w_stg_2_0_26, w_stg_2_1_26, w_stg_2_2_26);
	full_adder_md fa566( w_stg_3_5_26, w_stg_3_1_27, w_stg_2_3_26, w_stg_2_4_26, w_stg_2_5_26);
	full_adder_md fa567( w_stg_3_6_26, w_stg_3_2_27, w_stg_2_6_26, w_stg_2_7_26, w_stg_2_8_26);
	full_adder_md fa568( w_stg_3_7_26, w_stg_3_3_27, w_stg_2_9_26, w_stg_2_10_26, w_stg_2_11_26);
	full_adder_md fa569( w_stg_3_4_27, w_stg_3_0_28, w_stg_2_0_27, w_stg_2_1_27, w_stg_2_2_27);
	full_adder_md fa570( w_stg_3_5_27, w_stg_3_1_28, w_stg_2_3_27, w_stg_2_4_27, w_stg_2_5_27);
	full_adder_md fa571( w_stg_3_6_27, w_stg_3_2_28, w_stg_2_6_27, w_stg_2_7_27, w_stg_2_8_27);
	full_adder_md fa572( w_stg_3_7_27, w_stg_3_3_28, w_stg_2_9_27, w_stg_2_10_27, w_stg_2_11_27);
	assign w_stg_3_8_27 = w_stg_2_12_27;
	full_adder_md fa573( w_stg_3_4_28, w_stg_3_0_29, w_stg_2_0_28, w_stg_2_1_28, w_stg_2_2_28);
	full_adder_md fa574( w_stg_3_5_28, w_stg_3_1_29, w_stg_2_3_28, w_stg_2_4_28, w_stg_2_5_28);
	full_adder_md fa575( w_stg_3_6_28, w_stg_3_2_29, w_stg_2_6_28, w_stg_2_7_28, w_stg_2_8_28);
	full_adder_md fa576( w_stg_3_7_28, w_stg_3_3_29, w_stg_2_9_28, w_stg_2_10_28, w_stg_2_11_28);
	assign w_stg_3_8_28 = w_stg_2_12_28;
	full_adder_md fa577( w_stg_3_4_29, w_stg_3_0_30, w_stg_2_0_29, w_stg_2_1_29, w_stg_2_2_29);
	full_adder_md fa578( w_stg_3_5_29, w_stg_3_1_30, w_stg_2_3_29, w_stg_2_4_29, w_stg_2_5_29);
	full_adder_md fa579( w_stg_3_6_29, w_stg_3_2_30, w_stg_2_6_29, w_stg_2_7_29, w_stg_2_8_29);
	full_adder_md fa580( w_stg_3_7_29, w_stg_3_3_30, w_stg_2_9_29, w_stg_2_10_29, w_stg_2_11_29);
	assign w_stg_3_8_29 = w_stg_2_12_29;
	full_adder_md fa581( w_stg_3_4_30, w_stg_3_0_31, w_stg_2_0_30, w_stg_2_1_30, w_stg_2_2_30);
	full_adder_md fa582( w_stg_3_5_30, w_stg_3_1_31, w_stg_2_3_30, w_stg_2_4_30, w_stg_2_5_30);
	full_adder_md fa583( w_stg_3_6_30, w_stg_3_2_31, w_stg_2_6_30, w_stg_2_7_30, w_stg_2_8_30);
	full_adder_md fa584( w_stg_3_7_30, w_stg_3_3_31, w_stg_2_9_30, w_stg_2_10_30, w_stg_2_11_30);
	half_adder ha82( w_stg_3_8_30, w_stg_3_4_31, w_stg_2_12_30, w_stg_2_13_30);
	full_adder_md fa585( w_stg_3_5_31, w_stg_3_0_32, w_stg_2_0_31, w_stg_2_1_31, w_stg_2_2_31);
	full_adder_md fa586( w_stg_3_6_31, w_stg_3_1_32, w_stg_2_3_31, w_stg_2_4_31, w_stg_2_5_31);
	full_adder_md fa587( w_stg_3_7_31, w_stg_3_2_32, w_stg_2_6_31, w_stg_2_7_31, w_stg_2_8_31);
	full_adder_md fa588( w_stg_3_8_31, w_stg_3_3_32, w_stg_2_9_31, w_stg_2_10_31, w_stg_2_11_31);
	half_adder ha83( w_stg_3_9_31, w_stg_3_4_32, w_stg_2_12_31, w_stg_2_13_31);
	full_adder_md fa589( w_stg_3_5_32, w_stg_3_0_33, w_stg_2_0_32, w_stg_2_1_32, w_stg_2_2_32);
	full_adder_md fa590( w_stg_3_6_32, w_stg_3_1_33, w_stg_2_3_32, w_stg_2_4_32, w_stg_2_5_32);
	full_adder_md fa591( w_stg_3_7_32, w_stg_3_2_33, w_stg_2_6_32, w_stg_2_7_32, w_stg_2_8_32);
	full_adder_md fa592( w_stg_3_8_32, w_stg_3_3_33, w_stg_2_9_32, w_stg_2_10_32, w_stg_2_11_32);
	full_adder_md fa593( w_stg_3_9_32, w_stg_3_4_33, w_stg_2_12_32, w_stg_2_13_32, w_stg_2_14_32);
	full_adder_md fa594( w_stg_3_5_33, w_stg_3_0_34, w_stg_2_0_33, w_stg_2_1_33, w_stg_2_2_33);
	full_adder_md fa595( w_stg_3_6_33, w_stg_3_1_34, w_stg_2_3_33, w_stg_2_4_33, w_stg_2_5_33);
	full_adder_md fa596( w_stg_3_7_33, w_stg_3_2_34, w_stg_2_6_33, w_stg_2_7_33, w_stg_2_8_33);
	full_adder_md fa597( w_stg_3_8_33, w_stg_3_3_34, w_stg_2_9_33, w_stg_2_10_33, w_stg_2_11_33);
	full_adder_md fa598( w_stg_3_9_33, w_stg_3_4_34, w_stg_2_12_33, w_stg_2_13_33, w_stg_2_14_33);
	full_adder_md fa599( w_stg_3_5_34, w_stg_3_0_35, w_stg_2_0_34, w_stg_2_1_34, w_stg_2_2_34);
	full_adder_md fa600( w_stg_3_6_34, w_stg_3_1_35, w_stg_2_3_34, w_stg_2_4_34, w_stg_2_5_34);
	full_adder_md fa601( w_stg_3_7_34, w_stg_3_2_35, w_stg_2_6_34, w_stg_2_7_34, w_stg_2_8_34);
	full_adder_md fa602( w_stg_3_8_34, w_stg_3_3_35, w_stg_2_9_34, w_stg_2_10_34, w_stg_2_11_34);
	half_adder ha84( w_stg_3_9_34, w_stg_3_4_35, w_stg_2_12_34, w_stg_2_13_34);
	full_adder_md fa603( w_stg_3_5_35, w_stg_3_0_36, w_stg_2_0_35, w_stg_2_1_35, w_stg_2_2_35);
	full_adder_md fa604( w_stg_3_6_35, w_stg_3_1_36, w_stg_2_3_35, w_stg_2_4_35, w_stg_2_5_35);
	full_adder_md fa605( w_stg_3_7_35, w_stg_3_2_36, w_stg_2_6_35, w_stg_2_7_35, w_stg_2_8_35);
	full_adder_md fa606( w_stg_3_8_35, w_stg_3_3_36, w_stg_2_9_35, w_stg_2_10_35, w_stg_2_11_35);
	half_adder ha85( w_stg_3_9_35, w_stg_3_4_36, w_stg_2_12_35, w_stg_2_13_35);
	full_adder_md fa607( w_stg_3_5_36, w_stg_3_0_37, w_stg_2_0_36, w_stg_2_1_36, w_stg_2_2_36);
	full_adder_md fa608( w_stg_3_6_36, w_stg_3_1_37, w_stg_2_3_36, w_stg_2_4_36, w_stg_2_5_36);
	full_adder_md fa609( w_stg_3_7_36, w_stg_3_2_37, w_stg_2_6_36, w_stg_2_7_36, w_stg_2_8_36);
	full_adder_md fa610( w_stg_3_8_36, w_stg_3_3_37, w_stg_2_9_36, w_stg_2_10_36, w_stg_2_11_36);
	half_adder ha86( w_stg_3_9_36, w_stg_3_4_37, w_stg_2_12_36, w_stg_2_13_36);
	full_adder_md fa611( w_stg_3_5_37, w_stg_3_0_38, w_stg_2_0_37, w_stg_2_1_37, w_stg_2_2_37);
	full_adder_md fa612( w_stg_3_6_37, w_stg_3_1_38, w_stg_2_3_37, w_stg_2_4_37, w_stg_2_5_37);
	full_adder_md fa613( w_stg_3_7_37, w_stg_3_2_38, w_stg_2_6_37, w_stg_2_7_37, w_stg_2_8_37);
	full_adder_md fa614( w_stg_3_8_37, w_stg_3_3_38, w_stg_2_9_37, w_stg_2_10_37, w_stg_2_11_37);
	assign w_stg_3_9_37 = w_stg_2_12_37;
	full_adder_md fa615( w_stg_3_4_38, w_stg_3_0_39, w_stg_2_0_38, w_stg_2_1_38, w_stg_2_2_38);
	full_adder_md fa616( w_stg_3_5_38, w_stg_3_1_39, w_stg_2_3_38, w_stg_2_4_38, w_stg_2_5_38);
	full_adder_md fa617( w_stg_3_6_38, w_stg_3_2_39, w_stg_2_6_38, w_stg_2_7_38, w_stg_2_8_38);
	full_adder_md fa618( w_stg_3_7_38, w_stg_3_3_39, w_stg_2_9_38, w_stg_2_10_38, w_stg_2_11_38);
	full_adder_md fa619( w_stg_3_4_39, w_stg_3_0_40, w_stg_2_0_39, w_stg_2_1_39, w_stg_2_2_39);
	full_adder_md fa620( w_stg_3_5_39, w_stg_3_1_40, w_stg_2_3_39, w_stg_2_4_39, w_stg_2_5_39);
	full_adder_md fa621( w_stg_3_6_39, w_stg_3_2_40, w_stg_2_6_39, w_stg_2_7_39, w_stg_2_8_39);
	full_adder_md fa622( w_stg_3_7_39, w_stg_3_3_40, w_stg_2_9_39, w_stg_2_10_39, w_stg_2_11_39);
	full_adder_md fa623( w_stg_3_4_40, w_stg_3_0_41, w_stg_2_0_40, w_stg_2_1_40, w_stg_2_2_40);
	full_adder_md fa624( w_stg_3_5_40, w_stg_3_1_41, w_stg_2_3_40, w_stg_2_4_40, w_stg_2_5_40);
	full_adder_md fa625( w_stg_3_6_40, w_stg_3_2_41, w_stg_2_6_40, w_stg_2_7_40, w_stg_2_8_40);
	full_adder_md fa626( w_stg_3_7_40, w_stg_3_3_41, w_stg_2_9_40, w_stg_2_10_40, w_stg_2_11_40);
	full_adder_md fa627( w_stg_3_4_41, w_stg_3_0_42, w_stg_2_0_41, w_stg_2_1_41, w_stg_2_2_41);
	full_adder_md fa628( w_stg_3_5_41, w_stg_3_1_42, w_stg_2_3_41, w_stg_2_4_41, w_stg_2_5_41);
	full_adder_md fa629( w_stg_3_6_41, w_stg_3_2_42, w_stg_2_6_41, w_stg_2_7_41, w_stg_2_8_41);
	half_adder ha87( w_stg_3_7_41, w_stg_3_3_42, w_stg_2_9_41, w_stg_2_10_41);
	full_adder_md fa630( w_stg_3_4_42, w_stg_3_0_43, w_stg_2_0_42, w_stg_2_1_42, w_stg_2_2_42);
	full_adder_md fa631( w_stg_3_5_42, w_stg_3_1_43, w_stg_2_3_42, w_stg_2_4_42, w_stg_2_5_42);
	full_adder_md fa632( w_stg_3_6_42, w_stg_3_2_43, w_stg_2_6_42, w_stg_2_7_42, w_stg_2_8_42);
	half_adder ha88( w_stg_3_7_42, w_stg_3_3_43, w_stg_2_9_42, w_stg_2_10_42);
	full_adder_md fa633( w_stg_3_4_43, w_stg_3_0_44, w_stg_2_0_43, w_stg_2_1_43, w_stg_2_2_43);
	full_adder_md fa634( w_stg_3_5_43, w_stg_3_1_44, w_stg_2_3_43, w_stg_2_4_43, w_stg_2_5_43);
	full_adder_md fa635( w_stg_3_6_43, w_stg_3_2_44, w_stg_2_6_43, w_stg_2_7_43, w_stg_2_8_43);
	assign w_stg_3_7_43 = w_stg_2_9_43;
	full_adder_md fa636( w_stg_3_3_44, w_stg_3_0_45, w_stg_2_0_44, w_stg_2_1_44, w_stg_2_2_44);
	full_adder_md fa637( w_stg_3_4_44, w_stg_3_1_45, w_stg_2_3_44, w_stg_2_4_44, w_stg_2_5_44);
	full_adder_md fa638( w_stg_3_5_44, w_stg_3_2_45, w_stg_2_6_44, w_stg_2_7_44, w_stg_2_8_44);
	assign w_stg_3_6_44 = w_stg_2_9_44;
	full_adder_md fa639( w_stg_3_3_45, w_stg_3_0_46, w_stg_2_0_45, w_stg_2_1_45, w_stg_2_2_45);
	full_adder_md fa640( w_stg_3_4_45, w_stg_3_1_46, w_stg_2_3_45, w_stg_2_4_45, w_stg_2_5_45);
	full_adder_md fa641( w_stg_3_5_45, w_stg_3_2_46, w_stg_2_6_45, w_stg_2_7_45, w_stg_2_8_45);
	assign w_stg_3_6_45 = w_stg_2_9_45;
	full_adder_md fa642( w_stg_3_3_46, w_stg_3_0_47, w_stg_2_0_46, w_stg_2_1_46, w_stg_2_2_46);
	full_adder_md fa643( w_stg_3_4_46, w_stg_3_1_47, w_stg_2_3_46, w_stg_2_4_46, w_stg_2_5_46);
	full_adder_md fa644( w_stg_3_5_46, w_stg_3_2_47, w_stg_2_6_46, w_stg_2_7_46, w_stg_2_8_46);
	full_adder_md fa645( w_stg_3_3_47, w_stg_3_0_48, w_stg_2_0_47, w_stg_2_1_47, w_stg_2_2_47);
	full_adder_md fa646( w_stg_3_4_47, w_stg_3_1_48, w_stg_2_3_47, w_stg_2_4_47, w_stg_2_5_47);
	half_adder ha89( w_stg_3_5_47, w_stg_3_2_48, w_stg_2_6_47, w_stg_2_7_47);
	full_adder_md fa647( w_stg_3_3_48, w_stg_3_0_49, w_stg_2_0_48, w_stg_2_1_48, w_stg_2_2_48);
	full_adder_md fa648( w_stg_3_4_48, w_stg_3_1_49, w_stg_2_3_48, w_stg_2_4_48, w_stg_2_5_48);
	half_adder ha90( w_stg_3_5_48, w_stg_3_2_49, w_stg_2_6_48, w_stg_2_7_48);
	full_adder_md fa649( w_stg_3_3_49, w_stg_3_0_50, w_stg_2_0_49, w_stg_2_1_49, w_stg_2_2_49);
	full_adder_md fa650( w_stg_3_4_49, w_stg_3_1_50, w_stg_2_3_49, w_stg_2_4_49, w_stg_2_5_49);
	half_adder ha91( w_stg_3_5_49, w_stg_3_2_50, w_stg_2_6_49, w_stg_2_7_49);
	full_adder_md fa651( w_stg_3_3_50, w_stg_3_0_51, w_stg_2_0_50, w_stg_2_1_50, w_stg_2_2_50);
	full_adder_md fa652( w_stg_3_4_50, w_stg_3_1_51, w_stg_2_3_50, w_stg_2_4_50, w_stg_2_5_50);
	assign w_stg_3_5_50 = w_stg_2_6_50;
	full_adder_md fa653( w_stg_3_2_51, w_stg_3_0_52, w_stg_2_0_51, w_stg_2_1_51, w_stg_2_2_51);
	full_adder_md fa654( w_stg_3_3_51, w_stg_3_1_52, w_stg_2_3_51, w_stg_2_4_51, w_stg_2_5_51);
	assign w_stg_3_4_51 = w_stg_2_6_51;
	full_adder_md fa655( w_stg_3_2_52, w_stg_3_0_53, w_stg_2_0_52, w_stg_2_1_52, w_stg_2_2_52);
	full_adder_md fa656( w_stg_3_3_52, w_stg_3_1_53, w_stg_2_3_52, w_stg_2_4_52, w_stg_2_5_52);
	full_adder_md fa657( w_stg_3_2_53, w_stg_3_0_54, w_stg_2_0_53, w_stg_2_1_53, w_stg_2_2_53);
	full_adder_md fa658( w_stg_3_3_53, w_stg_3_1_54, w_stg_2_3_53, w_stg_2_4_53, w_stg_2_5_53);
	full_adder_md fa659( w_stg_3_2_54, w_stg_3_0_55, w_stg_2_0_54, w_stg_2_1_54, w_stg_2_2_54);
	full_adder_md fa660( w_stg_3_3_54, w_stg_3_1_55, w_stg_2_3_54, w_stg_2_4_54, w_stg_2_5_54);
	full_adder_md fa661( w_stg_3_2_55, w_stg_3_0_56, w_stg_2_0_55, w_stg_2_1_55, w_stg_2_2_55);
	half_adder ha92( w_stg_3_3_55, w_stg_3_1_56, w_stg_2_3_55, w_stg_2_4_55);
	full_adder_md fa662( w_stg_3_2_56, w_stg_3_0_57, w_stg_2_0_56, w_stg_2_1_56, w_stg_2_2_56);
	assign w_stg_3_3_56 = w_stg_2_3_56;
	full_adder_md fa663( w_stg_3_1_57, w_stg_3_0_58, w_stg_2_0_57, w_stg_2_1_57, w_stg_2_2_57);
	assign w_stg_3_2_57 = w_stg_2_3_57;
	full_adder_md fa664( w_stg_3_1_58, w_stg_3_0_59, w_stg_2_0_58, w_stg_2_1_58, w_stg_2_2_58);
	assign w_stg_3_2_58 = w_stg_2_3_58;
	full_adder_md fa665( w_stg_3_1_59, w_stg_3_0_60, w_stg_2_0_59, w_stg_2_1_59, w_stg_2_2_59);
	full_adder_md fa666( w_stg_3_1_60, w_stg_3_0_61, w_stg_2_0_60, w_stg_2_1_60, w_stg_2_2_60);
	half_adder ha93( w_stg_3_1_61, w_stg_3_0_62, w_stg_2_0_61, w_stg_2_1_61);
	half_adder ha94( w_stg_3_1_62, w_stg_3_0_63, w_stg_2_0_62, w_stg_2_1_62);
	assign w_stg_3_1_63 = w_stg_2_0_63;
	assign w_stg_4_0_0 = w_stg_3_0_0;
	assign w_stg_4_0_1 = w_stg_3_0_1;
	assign w_stg_4_0_2 = w_stg_3_0_2;
	assign w_stg_4_0_3 = w_stg_3_0_3;
	half_adder ha95( w_stg_4_0_4, w_stg_4_0_5, w_stg_3_0_4, w_stg_3_1_4);
	half_adder ha96( w_stg_4_1_5, w_stg_4_0_6, w_stg_3_0_5, w_stg_3_1_5);
	half_adder ha97( w_stg_4_1_6, w_stg_4_0_7, w_stg_3_0_6, w_stg_3_1_6);
	full_adder_md fa667( w_stg_4_1_7, w_stg_4_0_8, w_stg_3_0_7, w_stg_3_1_7, w_stg_3_2_7);
	full_adder_md fa668( w_stg_4_1_8, w_stg_4_0_9, w_stg_3_0_8, w_stg_3_1_8, w_stg_3_2_8);
	full_adder_md fa669( w_stg_4_1_9, w_stg_4_0_10, w_stg_3_0_9, w_stg_3_1_9, w_stg_3_2_9);
	full_adder_md fa670( w_stg_4_1_10, w_stg_4_0_11, w_stg_3_0_10, w_stg_3_1_10, w_stg_3_2_10);
	assign w_stg_4_2_10 = w_stg_3_3_10;
	full_adder_md fa671( w_stg_4_1_11, w_stg_4_0_12, w_stg_3_0_11, w_stg_3_1_11, w_stg_3_2_11);
	assign w_stg_4_2_11 = w_stg_3_3_11;
	full_adder_md fa672( w_stg_4_1_12, w_stg_4_0_13, w_stg_3_0_12, w_stg_3_1_12, w_stg_3_2_12);
	assign w_stg_4_2_12 = w_stg_3_3_12;
	full_adder_md fa673( w_stg_4_1_13, w_stg_4_0_14, w_stg_3_0_13, w_stg_3_1_13, w_stg_3_2_13);
	assign w_stg_4_2_13 = w_stg_3_3_13;
	full_adder_md fa674( w_stg_4_1_14, w_stg_4_0_15, w_stg_3_0_14, w_stg_3_1_14, w_stg_3_2_14);
	half_adder ha98( w_stg_4_2_14, w_stg_4_1_15, w_stg_3_3_14, w_stg_3_4_14);
	full_adder_md fa675( w_stg_4_2_15, w_stg_4_0_16, w_stg_3_0_15, w_stg_3_1_15, w_stg_3_2_15);
	half_adder ha99( w_stg_4_3_15, w_stg_4_1_16, w_stg_3_3_15, w_stg_3_4_15);
	full_adder_md fa676( w_stg_4_2_16, w_stg_4_0_17, w_stg_3_0_16, w_stg_3_1_16, w_stg_3_2_16);
	half_adder ha100( w_stg_4_3_16, w_stg_4_1_17, w_stg_3_3_16, w_stg_3_4_16);
	full_adder_md fa677( w_stg_4_2_17, w_stg_4_0_18, w_stg_3_0_17, w_stg_3_1_17, w_stg_3_2_17);
	full_adder_md fa678( w_stg_4_3_17, w_stg_4_1_18, w_stg_3_3_17, w_stg_3_4_17, w_stg_3_5_17);
	full_adder_md fa679( w_stg_4_2_18, w_stg_4_0_19, w_stg_3_0_18, w_stg_3_1_18, w_stg_3_2_18);
	full_adder_md fa680( w_stg_4_3_18, w_stg_4_1_19, w_stg_3_3_18, w_stg_3_4_18, w_stg_3_5_18);
	full_adder_md fa681( w_stg_4_2_19, w_stg_4_0_20, w_stg_3_0_19, w_stg_3_1_19, w_stg_3_2_19);
	full_adder_md fa682( w_stg_4_3_19, w_stg_4_1_20, w_stg_3_3_19, w_stg_3_4_19, w_stg_3_5_19);
	full_adder_md fa683( w_stg_4_2_20, w_stg_4_0_21, w_stg_3_0_20, w_stg_3_1_20, w_stg_3_2_20);
	full_adder_md fa684( w_stg_4_3_20, w_stg_4_1_21, w_stg_3_3_20, w_stg_3_4_20, w_stg_3_5_20);
	full_adder_md fa685( w_stg_4_2_21, w_stg_4_0_22, w_stg_3_0_21, w_stg_3_1_21, w_stg_3_2_21);
	full_adder_md fa686( w_stg_4_3_21, w_stg_4_1_22, w_stg_3_3_21, w_stg_3_4_21, w_stg_3_5_21);
	assign w_stg_4_4_21 = w_stg_3_6_21;
	full_adder_md fa687( w_stg_4_2_22, w_stg_4_0_23, w_stg_3_0_22, w_stg_3_1_22, w_stg_3_2_22);
	full_adder_md fa688( w_stg_4_3_22, w_stg_4_1_23, w_stg_3_3_22, w_stg_3_4_22, w_stg_3_5_22);
	assign w_stg_4_4_22 = w_stg_3_6_22;
	full_adder_md fa689( w_stg_4_2_23, w_stg_4_0_24, w_stg_3_0_23, w_stg_3_1_23, w_stg_3_2_23);
	full_adder_md fa690( w_stg_4_3_23, w_stg_4_1_24, w_stg_3_3_23, w_stg_3_4_23, w_stg_3_5_23);
	assign w_stg_4_4_23 = w_stg_3_6_23;
	full_adder_md fa691( w_stg_4_2_24, w_stg_4_0_25, w_stg_3_0_24, w_stg_3_1_24, w_stg_3_2_24);
	full_adder_md fa692( w_stg_4_3_24, w_stg_4_1_25, w_stg_3_3_24, w_stg_3_4_24, w_stg_3_5_24);
	half_adder ha101( w_stg_4_4_24, w_stg_4_2_25, w_stg_3_6_24, w_stg_3_7_24);
	full_adder_md fa693( w_stg_4_3_25, w_stg_4_0_26, w_stg_3_0_25, w_stg_3_1_25, w_stg_3_2_25);
	full_adder_md fa694( w_stg_4_4_25, w_stg_4_1_26, w_stg_3_3_25, w_stg_3_4_25, w_stg_3_5_25);
	half_adder ha102( w_stg_4_5_25, w_stg_4_2_26, w_stg_3_6_25, w_stg_3_7_25);
	full_adder_md fa695( w_stg_4_3_26, w_stg_4_0_27, w_stg_3_0_26, w_stg_3_1_26, w_stg_3_2_26);
	full_adder_md fa696( w_stg_4_4_26, w_stg_4_1_27, w_stg_3_3_26, w_stg_3_4_26, w_stg_3_5_26);
	half_adder ha103( w_stg_4_5_26, w_stg_4_2_27, w_stg_3_6_26, w_stg_3_7_26);
	full_adder_md fa697( w_stg_4_3_27, w_stg_4_0_28, w_stg_3_0_27, w_stg_3_1_27, w_stg_3_2_27);
	full_adder_md fa698( w_stg_4_4_27, w_stg_4_1_28, w_stg_3_3_27, w_stg_3_4_27, w_stg_3_5_27);
	full_adder_md fa699( w_stg_4_5_27, w_stg_4_2_28, w_stg_3_6_27, w_stg_3_7_27, w_stg_3_8_27);
	full_adder_md fa700( w_stg_4_3_28, w_stg_4_0_29, w_stg_3_0_28, w_stg_3_1_28, w_stg_3_2_28);
	full_adder_md fa701( w_stg_4_4_28, w_stg_4_1_29, w_stg_3_3_28, w_stg_3_4_28, w_stg_3_5_28);
	full_adder_md fa702( w_stg_4_5_28, w_stg_4_2_29, w_stg_3_6_28, w_stg_3_7_28, w_stg_3_8_28);
	full_adder_md fa703( w_stg_4_3_29, w_stg_4_0_30, w_stg_3_0_29, w_stg_3_1_29, w_stg_3_2_29);
	full_adder_md fa704( w_stg_4_4_29, w_stg_4_1_30, w_stg_3_3_29, w_stg_3_4_29, w_stg_3_5_29);
	full_adder_md fa705( w_stg_4_5_29, w_stg_4_2_30, w_stg_3_6_29, w_stg_3_7_29, w_stg_3_8_29);
	full_adder_md fa706( w_stg_4_3_30, w_stg_4_0_31, w_stg_3_0_30, w_stg_3_1_30, w_stg_3_2_30);
	full_adder_md fa707( w_stg_4_4_30, w_stg_4_1_31, w_stg_3_3_30, w_stg_3_4_30, w_stg_3_5_30);
	full_adder_md fa708( w_stg_4_5_30, w_stg_4_2_31, w_stg_3_6_30, w_stg_3_7_30, w_stg_3_8_30);
	full_adder_md fa709( w_stg_4_3_31, w_stg_4_0_32, w_stg_3_0_31, w_stg_3_1_31, w_stg_3_2_31);
	full_adder_md fa710( w_stg_4_4_31, w_stg_4_1_32, w_stg_3_3_31, w_stg_3_4_31, w_stg_3_5_31);
	full_adder_md fa711( w_stg_4_5_31, w_stg_4_2_32, w_stg_3_6_31, w_stg_3_7_31, w_stg_3_8_31);
	assign w_stg_4_6_31 = w_stg_3_9_31;
	full_adder_md fa712( w_stg_4_3_32, w_stg_4_0_33, w_stg_3_0_32, w_stg_3_1_32, w_stg_3_2_32);
	full_adder_md fa713( w_stg_4_4_32, w_stg_4_1_33, w_stg_3_3_32, w_stg_3_4_32, w_stg_3_5_32);
	full_adder_md fa714( w_stg_4_5_32, w_stg_4_2_33, w_stg_3_6_32, w_stg_3_7_32, w_stg_3_8_32);
	assign w_stg_4_6_32 = w_stg_3_9_32;
	full_adder_md fa715( w_stg_4_3_33, w_stg_4_0_34, w_stg_3_0_33, w_stg_3_1_33, w_stg_3_2_33);
	full_adder_md fa716( w_stg_4_4_33, w_stg_4_1_34, w_stg_3_3_33, w_stg_3_4_33, w_stg_3_5_33);
	full_adder_md fa717( w_stg_4_5_33, w_stg_4_2_34, w_stg_3_6_33, w_stg_3_7_33, w_stg_3_8_33);
	assign w_stg_4_6_33 = w_stg_3_9_33;
	full_adder_md fa718( w_stg_4_3_34, w_stg_4_0_35, w_stg_3_0_34, w_stg_3_1_34, w_stg_3_2_34);
	full_adder_md fa719( w_stg_4_4_34, w_stg_4_1_35, w_stg_3_3_34, w_stg_3_4_34, w_stg_3_5_34);
	full_adder_md fa720( w_stg_4_5_34, w_stg_4_2_35, w_stg_3_6_34, w_stg_3_7_34, w_stg_3_8_34);
	assign w_stg_4_6_34 = w_stg_3_9_34;
	full_adder_md fa721( w_stg_4_3_35, w_stg_4_0_36, w_stg_3_0_35, w_stg_3_1_35, w_stg_3_2_35);
	full_adder_md fa722( w_stg_4_4_35, w_stg_4_1_36, w_stg_3_3_35, w_stg_3_4_35, w_stg_3_5_35);
	full_adder_md fa723( w_stg_4_5_35, w_stg_4_2_36, w_stg_3_6_35, w_stg_3_7_35, w_stg_3_8_35);
	assign w_stg_4_6_35 = w_stg_3_9_35;
	full_adder_md fa724( w_stg_4_3_36, w_stg_4_0_37, w_stg_3_0_36, w_stg_3_1_36, w_stg_3_2_36);
	full_adder_md fa725( w_stg_4_4_36, w_stg_4_1_37, w_stg_3_3_36, w_stg_3_4_36, w_stg_3_5_36);
	full_adder_md fa726( w_stg_4_5_36, w_stg_4_2_37, w_stg_3_6_36, w_stg_3_7_36, w_stg_3_8_36);
	assign w_stg_4_6_36 = w_stg_3_9_36;
	full_adder_md fa727( w_stg_4_3_37, w_stg_4_0_38, w_stg_3_0_37, w_stg_3_1_37, w_stg_3_2_37);
	full_adder_md fa728( w_stg_4_4_37, w_stg_4_1_38, w_stg_3_3_37, w_stg_3_4_37, w_stg_3_5_37);
	full_adder_md fa729( w_stg_4_5_37, w_stg_4_2_38, w_stg_3_6_37, w_stg_3_7_37, w_stg_3_8_37);
	assign w_stg_4_6_37 = w_stg_3_9_37;
	full_adder_md fa730( w_stg_4_3_38, w_stg_4_0_39, w_stg_3_0_38, w_stg_3_1_38, w_stg_3_2_38);
	full_adder_md fa731( w_stg_4_4_38, w_stg_4_1_39, w_stg_3_3_38, w_stg_3_4_38, w_stg_3_5_38);
	half_adder ha104( w_stg_4_5_38, w_stg_4_2_39, w_stg_3_6_38, w_stg_3_7_38);
	full_adder_md fa732( w_stg_4_3_39, w_stg_4_0_40, w_stg_3_0_39, w_stg_3_1_39, w_stg_3_2_39);
	full_adder_md fa733( w_stg_4_4_39, w_stg_4_1_40, w_stg_3_3_39, w_stg_3_4_39, w_stg_3_5_39);
	half_adder ha105( w_stg_4_5_39, w_stg_4_2_40, w_stg_3_6_39, w_stg_3_7_39);
	full_adder_md fa734( w_stg_4_3_40, w_stg_4_0_41, w_stg_3_0_40, w_stg_3_1_40, w_stg_3_2_40);
	full_adder_md fa735( w_stg_4_4_40, w_stg_4_1_41, w_stg_3_3_40, w_stg_3_4_40, w_stg_3_5_40);
	half_adder ha106( w_stg_4_5_40, w_stg_4_2_41, w_stg_3_6_40, w_stg_3_7_40);
	full_adder_md fa736( w_stg_4_3_41, w_stg_4_0_42, w_stg_3_0_41, w_stg_3_1_41, w_stg_3_2_41);
	full_adder_md fa737( w_stg_4_4_41, w_stg_4_1_42, w_stg_3_3_41, w_stg_3_4_41, w_stg_3_5_41);
	half_adder ha107( w_stg_4_5_41, w_stg_4_2_42, w_stg_3_6_41, w_stg_3_7_41);
	full_adder_md fa738( w_stg_4_3_42, w_stg_4_0_43, w_stg_3_0_42, w_stg_3_1_42, w_stg_3_2_42);
	full_adder_md fa739( w_stg_4_4_42, w_stg_4_1_43, w_stg_3_3_42, w_stg_3_4_42, w_stg_3_5_42);
	half_adder ha108( w_stg_4_5_42, w_stg_4_2_43, w_stg_3_6_42, w_stg_3_7_42);
	full_adder_md fa740( w_stg_4_3_43, w_stg_4_0_44, w_stg_3_0_43, w_stg_3_1_43, w_stg_3_2_43);
	full_adder_md fa741( w_stg_4_4_43, w_stg_4_1_44, w_stg_3_3_43, w_stg_3_4_43, w_stg_3_5_43);
	half_adder ha109( w_stg_4_5_43, w_stg_4_2_44, w_stg_3_6_43, w_stg_3_7_43);
	full_adder_md fa742( w_stg_4_3_44, w_stg_4_0_45, w_stg_3_0_44, w_stg_3_1_44, w_stg_3_2_44);
	full_adder_md fa743( w_stg_4_4_44, w_stg_4_1_45, w_stg_3_3_44, w_stg_3_4_44, w_stg_3_5_44);
	assign w_stg_4_5_44 = w_stg_3_6_44;
	full_adder_md fa744( w_stg_4_2_45, w_stg_4_0_46, w_stg_3_0_45, w_stg_3_1_45, w_stg_3_2_45);
	full_adder_md fa745( w_stg_4_3_45, w_stg_4_1_46, w_stg_3_3_45, w_stg_3_4_45, w_stg_3_5_45);
	assign w_stg_4_4_45 = w_stg_3_6_45;
	full_adder_md fa746( w_stg_4_2_46, w_stg_4_0_47, w_stg_3_0_46, w_stg_3_1_46, w_stg_3_2_46);
	full_adder_md fa747( w_stg_4_3_46, w_stg_4_1_47, w_stg_3_3_46, w_stg_3_4_46, w_stg_3_5_46);
	full_adder_md fa748( w_stg_4_2_47, w_stg_4_0_48, w_stg_3_0_47, w_stg_3_1_47, w_stg_3_2_47);
	full_adder_md fa749( w_stg_4_3_47, w_stg_4_1_48, w_stg_3_3_47, w_stg_3_4_47, w_stg_3_5_47);
	full_adder_md fa750( w_stg_4_2_48, w_stg_4_0_49, w_stg_3_0_48, w_stg_3_1_48, w_stg_3_2_48);
	full_adder_md fa751( w_stg_4_3_48, w_stg_4_1_49, w_stg_3_3_48, w_stg_3_4_48, w_stg_3_5_48);
	full_adder_md fa752( w_stg_4_2_49, w_stg_4_0_50, w_stg_3_0_49, w_stg_3_1_49, w_stg_3_2_49);
	full_adder_md fa753( w_stg_4_3_49, w_stg_4_1_50, w_stg_3_3_49, w_stg_3_4_49, w_stg_3_5_49);
	full_adder_md fa754( w_stg_4_2_50, w_stg_4_0_51, w_stg_3_0_50, w_stg_3_1_50, w_stg_3_2_50);
	full_adder_md fa755( w_stg_4_3_50, w_stg_4_1_51, w_stg_3_3_50, w_stg_3_4_50, w_stg_3_5_50);
	full_adder_md fa756( w_stg_4_2_51, w_stg_4_0_52, w_stg_3_0_51, w_stg_3_1_51, w_stg_3_2_51);
	half_adder ha110( w_stg_4_3_51, w_stg_4_1_52, w_stg_3_3_51, w_stg_3_4_51);
	full_adder_md fa757( w_stg_4_2_52, w_stg_4_0_53, w_stg_3_0_52, w_stg_3_1_52, w_stg_3_2_52);
	assign w_stg_4_3_52 = w_stg_3_3_52;
	full_adder_md fa758( w_stg_4_1_53, w_stg_4_0_54, w_stg_3_0_53, w_stg_3_1_53, w_stg_3_2_53);
	assign w_stg_4_2_53 = w_stg_3_3_53;
	full_adder_md fa759( w_stg_4_1_54, w_stg_4_0_55, w_stg_3_0_54, w_stg_3_1_54, w_stg_3_2_54);
	assign w_stg_4_2_54 = w_stg_3_3_54;
	full_adder_md fa760( w_stg_4_1_55, w_stg_4_0_56, w_stg_3_0_55, w_stg_3_1_55, w_stg_3_2_55);
	assign w_stg_4_2_55 = w_stg_3_3_55;
	full_adder_md fa761( w_stg_4_1_56, w_stg_4_0_57, w_stg_3_0_56, w_stg_3_1_56, w_stg_3_2_56);
	assign w_stg_4_2_56 = w_stg_3_3_56;
	full_adder_md fa762( w_stg_4_1_57, w_stg_4_0_58, w_stg_3_0_57, w_stg_3_1_57, w_stg_3_2_57);
	full_adder_md fa763( w_stg_4_1_58, w_stg_4_0_59, w_stg_3_0_58, w_stg_3_1_58, w_stg_3_2_58);
	half_adder ha111( w_stg_4_1_59, w_stg_4_0_60, w_stg_3_0_59, w_stg_3_1_59);
	half_adder ha112( w_stg_4_1_60, w_stg_4_0_61, w_stg_3_0_60, w_stg_3_1_60);
	half_adder ha113( w_stg_4_1_61, w_stg_4_0_62, w_stg_3_0_61, w_stg_3_1_61);
	half_adder ha114( w_stg_4_1_62, w_stg_4_0_63, w_stg_3_0_62, w_stg_3_1_62);
	half_adder ha115( w_stg_4_1_63, w_stg_4_0_64, w_stg_3_0_63, w_stg_3_1_63);
	assign w_stg_5_0_0 = w_stg_4_0_0;
	assign w_stg_5_0_1 = w_stg_4_0_1;
	assign w_stg_5_0_2 = w_stg_4_0_2;
	assign w_stg_5_0_3 = w_stg_4_0_3;
	assign w_stg_5_0_4 = w_stg_4_0_4;
	half_adder ha116( w_stg_5_0_5, w_stg_5_0_6, w_stg_4_0_5, w_stg_4_1_5);
	half_adder ha117( w_stg_5_1_6, w_stg_5_0_7, w_stg_4_0_6, w_stg_4_1_6);
	half_adder ha118( w_stg_5_1_7, w_stg_5_0_8, w_stg_4_0_7, w_stg_4_1_7);
	half_adder ha119( w_stg_5_1_8, w_stg_5_0_9, w_stg_4_0_8, w_stg_4_1_8);
	half_adder ha120( w_stg_5_1_9, w_stg_5_0_10, w_stg_4_0_9, w_stg_4_1_9);
	full_adder_md fa764( w_stg_5_1_10, w_stg_5_0_11, w_stg_4_0_10, w_stg_4_1_10, w_stg_4_2_10);
	full_adder_md fa765( w_stg_5_1_11, w_stg_5_0_12, w_stg_4_0_11, w_stg_4_1_11, w_stg_4_2_11);
	full_adder_md fa766( w_stg_5_1_12, w_stg_5_0_13, w_stg_4_0_12, w_stg_4_1_12, w_stg_4_2_12);
	full_adder_md fa767( w_stg_5_1_13, w_stg_5_0_14, w_stg_4_0_13, w_stg_4_1_13, w_stg_4_2_13);
	full_adder_md fa768( w_stg_5_1_14, w_stg_5_0_15, w_stg_4_0_14, w_stg_4_1_14, w_stg_4_2_14);
	full_adder_md fa769( w_stg_5_1_15, w_stg_5_0_16, w_stg_4_0_15, w_stg_4_1_15, w_stg_4_2_15);
	assign w_stg_5_2_15 = w_stg_4_3_15;
	full_adder_md fa770( w_stg_5_1_16, w_stg_5_0_17, w_stg_4_0_16, w_stg_4_1_16, w_stg_4_2_16);
	assign w_stg_5_2_16 = w_stg_4_3_16;
	full_adder_md fa771( w_stg_5_1_17, w_stg_5_0_18, w_stg_4_0_17, w_stg_4_1_17, w_stg_4_2_17);
	assign w_stg_5_2_17 = w_stg_4_3_17;
	full_adder_md fa772( w_stg_5_1_18, w_stg_5_0_19, w_stg_4_0_18, w_stg_4_1_18, w_stg_4_2_18);
	assign w_stg_5_2_18 = w_stg_4_3_18;
	full_adder_md fa773( w_stg_5_1_19, w_stg_5_0_20, w_stg_4_0_19, w_stg_4_1_19, w_stg_4_2_19);
	assign w_stg_5_2_19 = w_stg_4_3_19;
	full_adder_md fa774( w_stg_5_1_20, w_stg_5_0_21, w_stg_4_0_20, w_stg_4_1_20, w_stg_4_2_20);
	assign w_stg_5_2_20 = w_stg_4_3_20;
	full_adder_md fa775( w_stg_5_1_21, w_stg_5_0_22, w_stg_4_0_21, w_stg_4_1_21, w_stg_4_2_21);
	half_adder ha121( w_stg_5_2_21, w_stg_5_1_22, w_stg_4_3_21, w_stg_4_4_21);
	full_adder_md fa776( w_stg_5_2_22, w_stg_5_0_23, w_stg_4_0_22, w_stg_4_1_22, w_stg_4_2_22);
	half_adder ha122( w_stg_5_3_22, w_stg_5_1_23, w_stg_4_3_22, w_stg_4_4_22);
	full_adder_md fa777( w_stg_5_2_23, w_stg_5_0_24, w_stg_4_0_23, w_stg_4_1_23, w_stg_4_2_23);
	half_adder ha123( w_stg_5_3_23, w_stg_5_1_24, w_stg_4_3_23, w_stg_4_4_23);
	full_adder_md fa778( w_stg_5_2_24, w_stg_5_0_25, w_stg_4_0_24, w_stg_4_1_24, w_stg_4_2_24);
	half_adder ha124( w_stg_5_3_24, w_stg_5_1_25, w_stg_4_3_24, w_stg_4_4_24);
	full_adder_md fa779( w_stg_5_2_25, w_stg_5_0_26, w_stg_4_0_25, w_stg_4_1_25, w_stg_4_2_25);
	full_adder_md fa780( w_stg_5_3_25, w_stg_5_1_26, w_stg_4_3_25, w_stg_4_4_25, w_stg_4_5_25);
	full_adder_md fa781( w_stg_5_2_26, w_stg_5_0_27, w_stg_4_0_26, w_stg_4_1_26, w_stg_4_2_26);
	full_adder_md fa782( w_stg_5_3_26, w_stg_5_1_27, w_stg_4_3_26, w_stg_4_4_26, w_stg_4_5_26);
	full_adder_md fa783( w_stg_5_2_27, w_stg_5_0_28, w_stg_4_0_27, w_stg_4_1_27, w_stg_4_2_27);
	full_adder_md fa784( w_stg_5_3_27, w_stg_5_1_28, w_stg_4_3_27, w_stg_4_4_27, w_stg_4_5_27);
	full_adder_md fa785( w_stg_5_2_28, w_stg_5_0_29, w_stg_4_0_28, w_stg_4_1_28, w_stg_4_2_28);
	full_adder_md fa786( w_stg_5_3_28, w_stg_5_1_29, w_stg_4_3_28, w_stg_4_4_28, w_stg_4_5_28);
	full_adder_md fa787( w_stg_5_2_29, w_stg_5_0_30, w_stg_4_0_29, w_stg_4_1_29, w_stg_4_2_29);
	full_adder_md fa788( w_stg_5_3_29, w_stg_5_1_30, w_stg_4_3_29, w_stg_4_4_29, w_stg_4_5_29);
	full_adder_md fa789( w_stg_5_2_30, w_stg_5_0_31, w_stg_4_0_30, w_stg_4_1_30, w_stg_4_2_30);
	full_adder_md fa790( w_stg_5_3_30, w_stg_5_1_31, w_stg_4_3_30, w_stg_4_4_30, w_stg_4_5_30);
	full_adder_md fa791( w_stg_5_2_31, w_stg_5_0_32, w_stg_4_0_31, w_stg_4_1_31, w_stg_4_2_31);
	full_adder_md fa792( w_stg_5_3_31, w_stg_5_1_32, w_stg_4_3_31, w_stg_4_4_31, w_stg_4_5_31);
	assign w_stg_5_4_31 = w_stg_4_6_31;
	full_adder_md fa793( w_stg_5_2_32, w_stg_5_0_33, w_stg_4_0_32, w_stg_4_1_32, w_stg_4_2_32);
	full_adder_md fa794( w_stg_5_3_32, w_stg_5_1_33, w_stg_4_3_32, w_stg_4_4_32, w_stg_4_5_32);
	assign w_stg_5_4_32 = w_stg_4_6_32;
	full_adder_md fa795( w_stg_5_2_33, w_stg_5_0_34, w_stg_4_0_33, w_stg_4_1_33, w_stg_4_2_33);
	full_adder_md fa796( w_stg_5_3_33, w_stg_5_1_34, w_stg_4_3_33, w_stg_4_4_33, w_stg_4_5_33);
	assign w_stg_5_4_33 = w_stg_4_6_33;
	full_adder_md fa797( w_stg_5_2_34, w_stg_5_0_35, w_stg_4_0_34, w_stg_4_1_34, w_stg_4_2_34);
	full_adder_md fa798( w_stg_5_3_34, w_stg_5_1_35, w_stg_4_3_34, w_stg_4_4_34, w_stg_4_5_34);
	assign w_stg_5_4_34 = w_stg_4_6_34;
	full_adder_md fa799( w_stg_5_2_35, w_stg_5_0_36, w_stg_4_0_35, w_stg_4_1_35, w_stg_4_2_35);
	full_adder_md fa800( w_stg_5_3_35, w_stg_5_1_36, w_stg_4_3_35, w_stg_4_4_35, w_stg_4_5_35);
	assign w_stg_5_4_35 = w_stg_4_6_35;
	full_adder_md fa801( w_stg_5_2_36, w_stg_5_0_37, w_stg_4_0_36, w_stg_4_1_36, w_stg_4_2_36);
	full_adder_md fa802( w_stg_5_3_36, w_stg_5_1_37, w_stg_4_3_36, w_stg_4_4_36, w_stg_4_5_36);
	assign w_stg_5_4_36 = w_stg_4_6_36;
	full_adder_md fa803( w_stg_5_2_37, w_stg_5_0_38, w_stg_4_0_37, w_stg_4_1_37, w_stg_4_2_37);
	full_adder_md fa804( w_stg_5_3_37, w_stg_5_1_38, w_stg_4_3_37, w_stg_4_4_37, w_stg_4_5_37);
	assign w_stg_5_4_37 = w_stg_4_6_37;
	full_adder_md fa805( w_stg_5_2_38, w_stg_5_0_39, w_stg_4_0_38, w_stg_4_1_38, w_stg_4_2_38);
	full_adder_md fa806( w_stg_5_3_38, w_stg_5_1_39, w_stg_4_3_38, w_stg_4_4_38, w_stg_4_5_38);
	full_adder_md fa807( w_stg_5_2_39, w_stg_5_0_40, w_stg_4_0_39, w_stg_4_1_39, w_stg_4_2_39);
	full_adder_md fa808( w_stg_5_3_39, w_stg_5_1_40, w_stg_4_3_39, w_stg_4_4_39, w_stg_4_5_39);
	full_adder_md fa809( w_stg_5_2_40, w_stg_5_0_41, w_stg_4_0_40, w_stg_4_1_40, w_stg_4_2_40);
	full_adder_md fa810( w_stg_5_3_40, w_stg_5_1_41, w_stg_4_3_40, w_stg_4_4_40, w_stg_4_5_40);
	full_adder_md fa811( w_stg_5_2_41, w_stg_5_0_42, w_stg_4_0_41, w_stg_4_1_41, w_stg_4_2_41);
	full_adder_md fa812( w_stg_5_3_41, w_stg_5_1_42, w_stg_4_3_41, w_stg_4_4_41, w_stg_4_5_41);
	full_adder_md fa813( w_stg_5_2_42, w_stg_5_0_43, w_stg_4_0_42, w_stg_4_1_42, w_stg_4_2_42);
	full_adder_md fa814( w_stg_5_3_42, w_stg_5_1_43, w_stg_4_3_42, w_stg_4_4_42, w_stg_4_5_42);
	full_adder_md fa815( w_stg_5_2_43, w_stg_5_0_44, w_stg_4_0_43, w_stg_4_1_43, w_stg_4_2_43);
	full_adder_md fa816( w_stg_5_3_43, w_stg_5_1_44, w_stg_4_3_43, w_stg_4_4_43, w_stg_4_5_43);
	full_adder_md fa817( w_stg_5_2_44, w_stg_5_0_45, w_stg_4_0_44, w_stg_4_1_44, w_stg_4_2_44);
	full_adder_md fa818( w_stg_5_3_44, w_stg_5_1_45, w_stg_4_3_44, w_stg_4_4_44, w_stg_4_5_44);
	full_adder_md fa819( w_stg_5_2_45, w_stg_5_0_46, w_stg_4_0_45, w_stg_4_1_45, w_stg_4_2_45);
	half_adder ha125( w_stg_5_3_45, w_stg_5_1_46, w_stg_4_3_45, w_stg_4_4_45);
	full_adder_md fa820( w_stg_5_2_46, w_stg_5_0_47, w_stg_4_0_46, w_stg_4_1_46, w_stg_4_2_46);
	assign w_stg_5_3_46 = w_stg_4_3_46;
	full_adder_md fa821( w_stg_5_1_47, w_stg_5_0_48, w_stg_4_0_47, w_stg_4_1_47, w_stg_4_2_47);
	assign w_stg_5_2_47 = w_stg_4_3_47;
	full_adder_md fa822( w_stg_5_1_48, w_stg_5_0_49, w_stg_4_0_48, w_stg_4_1_48, w_stg_4_2_48);
	assign w_stg_5_2_48 = w_stg_4_3_48;
	full_adder_md fa823( w_stg_5_1_49, w_stg_5_0_50, w_stg_4_0_49, w_stg_4_1_49, w_stg_4_2_49);
	assign w_stg_5_2_49 = w_stg_4_3_49;
	full_adder_md fa824( w_stg_5_1_50, w_stg_5_0_51, w_stg_4_0_50, w_stg_4_1_50, w_stg_4_2_50);
	assign w_stg_5_2_50 = w_stg_4_3_50;
	full_adder_md fa825( w_stg_5_1_51, w_stg_5_0_52, w_stg_4_0_51, w_stg_4_1_51, w_stg_4_2_51);
	assign w_stg_5_2_51 = w_stg_4_3_51;
	full_adder_md fa826( w_stg_5_1_52, w_stg_5_0_53, w_stg_4_0_52, w_stg_4_1_52, w_stg_4_2_52);
	assign w_stg_5_2_52 = w_stg_4_3_52;
	full_adder_md fa827( w_stg_5_1_53, w_stg_5_0_54, w_stg_4_0_53, w_stg_4_1_53, w_stg_4_2_53);
	full_adder_md fa828( w_stg_5_1_54, w_stg_5_0_55, w_stg_4_0_54, w_stg_4_1_54, w_stg_4_2_54);
	full_adder_md fa829( w_stg_5_1_55, w_stg_5_0_56, w_stg_4_0_55, w_stg_4_1_55, w_stg_4_2_55);
	full_adder_md fa830( w_stg_5_1_56, w_stg_5_0_57, w_stg_4_0_56, w_stg_4_1_56, w_stg_4_2_56);
	half_adder ha126( w_stg_5_1_57, w_stg_5_0_58, w_stg_4_0_57, w_stg_4_1_57);
	half_adder ha127( w_stg_5_1_58, w_stg_5_0_59, w_stg_4_0_58, w_stg_4_1_58);
	half_adder ha128( w_stg_5_1_59, w_stg_5_0_60, w_stg_4_0_59, w_stg_4_1_59);
	half_adder ha129( w_stg_5_1_60, w_stg_5_0_61, w_stg_4_0_60, w_stg_4_1_60);
	half_adder ha130( w_stg_5_1_61, w_stg_5_0_62, w_stg_4_0_61, w_stg_4_1_61);
	half_adder ha131( w_stg_5_1_62, w_stg_5_0_63, w_stg_4_0_62, w_stg_4_1_62);
	half_adder ha132( w_stg_5_1_63, w_stg_5_0_64, w_stg_4_0_63, w_stg_4_1_63);
	assign w_stg_5_1_64 = w_stg_4_0_64;
	assign w_stg_6_0_0 = w_stg_5_0_0;
	assign w_stg_6_0_1 = w_stg_5_0_1;
	assign w_stg_6_0_2 = w_stg_5_0_2;
	assign w_stg_6_0_3 = w_stg_5_0_3;
	assign w_stg_6_0_4 = w_stg_5_0_4;
	assign w_stg_6_0_5 = w_stg_5_0_5;
	half_adder ha133( w_stg_6_0_6, w_stg_6_0_7, w_stg_5_0_6, w_stg_5_1_6);
	half_adder ha134( w_stg_6_1_7, w_stg_6_0_8, w_stg_5_0_7, w_stg_5_1_7);
	half_adder ha135( w_stg_6_1_8, w_stg_6_0_9, w_stg_5_0_8, w_stg_5_1_8);
	half_adder ha136( w_stg_6_1_9, w_stg_6_0_10, w_stg_5_0_9, w_stg_5_1_9);
	half_adder ha137( w_stg_6_1_10, w_stg_6_0_11, w_stg_5_0_10, w_stg_5_1_10);
	half_adder ha138( w_stg_6_1_11, w_stg_6_0_12, w_stg_5_0_11, w_stg_5_1_11);
	half_adder ha139( w_stg_6_1_12, w_stg_6_0_13, w_stg_5_0_12, w_stg_5_1_12);
	half_adder ha140( w_stg_6_1_13, w_stg_6_0_14, w_stg_5_0_13, w_stg_5_1_13);
	half_adder ha141( w_stg_6_1_14, w_stg_6_0_15, w_stg_5_0_14, w_stg_5_1_14);
	full_adder_md fa831( w_stg_6_1_15, w_stg_6_0_16, w_stg_5_0_15, w_stg_5_1_15, w_stg_5_2_15);
	full_adder_md fa832( w_stg_6_1_16, w_stg_6_0_17, w_stg_5_0_16, w_stg_5_1_16, w_stg_5_2_16);
	full_adder_md fa833( w_stg_6_1_17, w_stg_6_0_18, w_stg_5_0_17, w_stg_5_1_17, w_stg_5_2_17);
	full_adder_md fa834( w_stg_6_1_18, w_stg_6_0_19, w_stg_5_0_18, w_stg_5_1_18, w_stg_5_2_18);
	full_adder_md fa835( w_stg_6_1_19, w_stg_6_0_20, w_stg_5_0_19, w_stg_5_1_19, w_stg_5_2_19);
	full_adder_md fa836( w_stg_6_1_20, w_stg_6_0_21, w_stg_5_0_20, w_stg_5_1_20, w_stg_5_2_20);
	full_adder_md fa837( w_stg_6_1_21, w_stg_6_0_22, w_stg_5_0_21, w_stg_5_1_21, w_stg_5_2_21);
	full_adder_md fa838( w_stg_6_1_22, w_stg_6_0_23, w_stg_5_0_22, w_stg_5_1_22, w_stg_5_2_22);
	assign w_stg_6_2_22 = w_stg_5_3_22;
	full_adder_md fa839( w_stg_6_1_23, w_stg_6_0_24, w_stg_5_0_23, w_stg_5_1_23, w_stg_5_2_23);
	assign w_stg_6_2_23 = w_stg_5_3_23;
	full_adder_md fa840( w_stg_6_1_24, w_stg_6_0_25, w_stg_5_0_24, w_stg_5_1_24, w_stg_5_2_24);
	assign w_stg_6_2_24 = w_stg_5_3_24;
	full_adder_md fa841( w_stg_6_1_25, w_stg_6_0_26, w_stg_5_0_25, w_stg_5_1_25, w_stg_5_2_25);
	assign w_stg_6_2_25 = w_stg_5_3_25;
	full_adder_md fa842( w_stg_6_1_26, w_stg_6_0_27, w_stg_5_0_26, w_stg_5_1_26, w_stg_5_2_26);
	assign w_stg_6_2_26 = w_stg_5_3_26;
	full_adder_md fa843( w_stg_6_1_27, w_stg_6_0_28, w_stg_5_0_27, w_stg_5_1_27, w_stg_5_2_27);
	assign w_stg_6_2_27 = w_stg_5_3_27;
	full_adder_md fa844( w_stg_6_1_28, w_stg_6_0_29, w_stg_5_0_28, w_stg_5_1_28, w_stg_5_2_28);
	assign w_stg_6_2_28 = w_stg_5_3_28;
	full_adder_md fa845( w_stg_6_1_29, w_stg_6_0_30, w_stg_5_0_29, w_stg_5_1_29, w_stg_5_2_29);
	assign w_stg_6_2_29 = w_stg_5_3_29;
	full_adder_md fa846( w_stg_6_1_30, w_stg_6_0_31, w_stg_5_0_30, w_stg_5_1_30, w_stg_5_2_30);
	assign w_stg_6_2_30 = w_stg_5_3_30;
	full_adder_md fa847( w_stg_6_1_31, w_stg_6_0_32, w_stg_5_0_31, w_stg_5_1_31, w_stg_5_2_31);
	half_adder ha142( w_stg_6_2_31, w_stg_6_1_32, w_stg_5_3_31, w_stg_5_4_31);
	full_adder_md fa848( w_stg_6_2_32, w_stg_6_0_33, w_stg_5_0_32, w_stg_5_1_32, w_stg_5_2_32);
	half_adder ha143( w_stg_6_3_32, w_stg_6_1_33, w_stg_5_3_32, w_stg_5_4_32);
	full_adder_md fa849( w_stg_6_2_33, w_stg_6_0_34, w_stg_5_0_33, w_stg_5_1_33, w_stg_5_2_33);
	half_adder ha144( w_stg_6_3_33, w_stg_6_1_34, w_stg_5_3_33, w_stg_5_4_33);
	full_adder_md fa850( w_stg_6_2_34, w_stg_6_0_35, w_stg_5_0_34, w_stg_5_1_34, w_stg_5_2_34);
	half_adder ha145( w_stg_6_3_34, w_stg_6_1_35, w_stg_5_3_34, w_stg_5_4_34);
	full_adder_md fa851( w_stg_6_2_35, w_stg_6_0_36, w_stg_5_0_35, w_stg_5_1_35, w_stg_5_2_35);
	half_adder ha146( w_stg_6_3_35, w_stg_6_1_36, w_stg_5_3_35, w_stg_5_4_35);
	full_adder_md fa852( w_stg_6_2_36, w_stg_6_0_37, w_stg_5_0_36, w_stg_5_1_36, w_stg_5_2_36);
	half_adder ha147( w_stg_6_3_36, w_stg_6_1_37, w_stg_5_3_36, w_stg_5_4_36);
	full_adder_md fa853( w_stg_6_2_37, w_stg_6_0_38, w_stg_5_0_37, w_stg_5_1_37, w_stg_5_2_37);
	half_adder ha148( w_stg_6_3_37, w_stg_6_1_38, w_stg_5_3_37, w_stg_5_4_37);
	full_adder_md fa854( w_stg_6_2_38, w_stg_6_0_39, w_stg_5_0_38, w_stg_5_1_38, w_stg_5_2_38);
	assign w_stg_6_3_38 = w_stg_5_3_38;
	full_adder_md fa855( w_stg_6_1_39, w_stg_6_0_40, w_stg_5_0_39, w_stg_5_1_39, w_stg_5_2_39);
	assign w_stg_6_2_39 = w_stg_5_3_39;
	full_adder_md fa856( w_stg_6_1_40, w_stg_6_0_41, w_stg_5_0_40, w_stg_5_1_40, w_stg_5_2_40);
	assign w_stg_6_2_40 = w_stg_5_3_40;
	full_adder_md fa857( w_stg_6_1_41, w_stg_6_0_42, w_stg_5_0_41, w_stg_5_1_41, w_stg_5_2_41);
	assign w_stg_6_2_41 = w_stg_5_3_41;
	full_adder_md fa858( w_stg_6_1_42, w_stg_6_0_43, w_stg_5_0_42, w_stg_5_1_42, w_stg_5_2_42);
	assign w_stg_6_2_42 = w_stg_5_3_42;
	full_adder_md fa859( w_stg_6_1_43, w_stg_6_0_44, w_stg_5_0_43, w_stg_5_1_43, w_stg_5_2_43);
	assign w_stg_6_2_43 = w_stg_5_3_43;
	full_adder_md fa860( w_stg_6_1_44, w_stg_6_0_45, w_stg_5_0_44, w_stg_5_1_44, w_stg_5_2_44);
	assign w_stg_6_2_44 = w_stg_5_3_44;
	full_adder_md fa861( w_stg_6_1_45, w_stg_6_0_46, w_stg_5_0_45, w_stg_5_1_45, w_stg_5_2_45);
	assign w_stg_6_2_45 = w_stg_5_3_45;
	full_adder_md fa862( w_stg_6_1_46, w_stg_6_0_47, w_stg_5_0_46, w_stg_5_1_46, w_stg_5_2_46);
	assign w_stg_6_2_46 = w_stg_5_3_46;
	full_adder_md fa863( w_stg_6_1_47, w_stg_6_0_48, w_stg_5_0_47, w_stg_5_1_47, w_stg_5_2_47);
	full_adder_md fa864( w_stg_6_1_48, w_stg_6_0_49, w_stg_5_0_48, w_stg_5_1_48, w_stg_5_2_48);
	full_adder_md fa865( w_stg_6_1_49, w_stg_6_0_50, w_stg_5_0_49, w_stg_5_1_49, w_stg_5_2_49);
	full_adder_md fa866( w_stg_6_1_50, w_stg_6_0_51, w_stg_5_0_50, w_stg_5_1_50, w_stg_5_2_50);
	full_adder_md fa867( w_stg_6_1_51, w_stg_6_0_52, w_stg_5_0_51, w_stg_5_1_51, w_stg_5_2_51);
	full_adder_md fa868( w_stg_6_1_52, w_stg_6_0_53, w_stg_5_0_52, w_stg_5_1_52, w_stg_5_2_52);
	half_adder ha149( w_stg_6_1_53, w_stg_6_0_54, w_stg_5_0_53, w_stg_5_1_53);
	half_adder ha150( w_stg_6_1_54, w_stg_6_0_55, w_stg_5_0_54, w_stg_5_1_54);
	half_adder ha151( w_stg_6_1_55, w_stg_6_0_56, w_stg_5_0_55, w_stg_5_1_55);
	half_adder ha152( w_stg_6_1_56, w_stg_6_0_57, w_stg_5_0_56, w_stg_5_1_56);
	half_adder ha153( w_stg_6_1_57, w_stg_6_0_58, w_stg_5_0_57, w_stg_5_1_57);
	half_adder ha154( w_stg_6_1_58, w_stg_6_0_59, w_stg_5_0_58, w_stg_5_1_58);
	half_adder ha155( w_stg_6_1_59, w_stg_6_0_60, w_stg_5_0_59, w_stg_5_1_59);
	half_adder ha156( w_stg_6_1_60, w_stg_6_0_61, w_stg_5_0_60, w_stg_5_1_60);
	half_adder ha157( w_stg_6_1_61, w_stg_6_0_62, w_stg_5_0_61, w_stg_5_1_61);
	half_adder ha158( w_stg_6_1_62, w_stg_6_0_63, w_stg_5_0_62, w_stg_5_1_62);
	half_adder ha159( w_stg_6_1_63, w_stg_6_0_64, w_stg_5_0_63, w_stg_5_1_63);
	half_adder ha160( w_stg_6_1_64, w_stg_6_0_65, w_stg_5_0_64, w_stg_5_1_64);
	assign w_stg_7_0_0 = w_stg_6_0_0;
	assign w_stg_7_0_1 = w_stg_6_0_1;
	assign w_stg_7_0_2 = w_stg_6_0_2;
	assign w_stg_7_0_3 = w_stg_6_0_3;
	assign w_stg_7_0_4 = w_stg_6_0_4;
	assign w_stg_7_0_5 = w_stg_6_0_5;
	assign w_stg_7_0_6 = w_stg_6_0_6;
	half_adder ha161( w_stg_7_0_7, w_stg_7_0_8, w_stg_6_0_7, w_stg_6_1_7);
	half_adder ha162( w_stg_7_1_8, w_stg_7_0_9, w_stg_6_0_8, w_stg_6_1_8);
	half_adder ha163( w_stg_7_1_9, w_stg_7_0_10, w_stg_6_0_9, w_stg_6_1_9);
	half_adder ha164( w_stg_7_1_10, w_stg_7_0_11, w_stg_6_0_10, w_stg_6_1_10);
	half_adder ha165( w_stg_7_1_11, w_stg_7_0_12, w_stg_6_0_11, w_stg_6_1_11);
	half_adder ha166( w_stg_7_1_12, w_stg_7_0_13, w_stg_6_0_12, w_stg_6_1_12);
	half_adder ha167( w_stg_7_1_13, w_stg_7_0_14, w_stg_6_0_13, w_stg_6_1_13);
	half_adder ha168( w_stg_7_1_14, w_stg_7_0_15, w_stg_6_0_14, w_stg_6_1_14);
	half_adder ha169( w_stg_7_1_15, w_stg_7_0_16, w_stg_6_0_15, w_stg_6_1_15);
	half_adder ha170( w_stg_7_1_16, w_stg_7_0_17, w_stg_6_0_16, w_stg_6_1_16);
	half_adder ha171( w_stg_7_1_17, w_stg_7_0_18, w_stg_6_0_17, w_stg_6_1_17);
	half_adder ha172( w_stg_7_1_18, w_stg_7_0_19, w_stg_6_0_18, w_stg_6_1_18);
	half_adder ha173( w_stg_7_1_19, w_stg_7_0_20, w_stg_6_0_19, w_stg_6_1_19);
	half_adder ha174( w_stg_7_1_20, w_stg_7_0_21, w_stg_6_0_20, w_stg_6_1_20);
	half_adder ha175( w_stg_7_1_21, w_stg_7_0_22, w_stg_6_0_21, w_stg_6_1_21);
	full_adder_md fa869( w_stg_7_1_22, w_stg_7_0_23, w_stg_6_0_22, w_stg_6_1_22, w_stg_6_2_22);
	full_adder_md fa870( w_stg_7_1_23, w_stg_7_0_24, w_stg_6_0_23, w_stg_6_1_23, w_stg_6_2_23);
	full_adder_md fa871( w_stg_7_1_24, w_stg_7_0_25, w_stg_6_0_24, w_stg_6_1_24, w_stg_6_2_24);
	full_adder_md fa872( w_stg_7_1_25, w_stg_7_0_26, w_stg_6_0_25, w_stg_6_1_25, w_stg_6_2_25);
	full_adder_md fa873( w_stg_7_1_26, w_stg_7_0_27, w_stg_6_0_26, w_stg_6_1_26, w_stg_6_2_26);
	full_adder_md fa874( w_stg_7_1_27, w_stg_7_0_28, w_stg_6_0_27, w_stg_6_1_27, w_stg_6_2_27);
	full_adder_md fa875( w_stg_7_1_28, w_stg_7_0_29, w_stg_6_0_28, w_stg_6_1_28, w_stg_6_2_28);
	full_adder_md fa876( w_stg_7_1_29, w_stg_7_0_30, w_stg_6_0_29, w_stg_6_1_29, w_stg_6_2_29);
	full_adder_md fa877( w_stg_7_1_30, w_stg_7_0_31, w_stg_6_0_30, w_stg_6_1_30, w_stg_6_2_30);
	full_adder_md fa878( w_stg_7_1_31, w_stg_7_0_32, w_stg_6_0_31, w_stg_6_1_31, w_stg_6_2_31);
	full_adder_md fa879( w_stg_7_1_32, w_stg_7_0_33, w_stg_6_0_32, w_stg_6_1_32, w_stg_6_2_32);
	assign w_stg_7_2_32 = w_stg_6_3_32;
	full_adder_md fa880( w_stg_7_1_33, w_stg_7_0_34, w_stg_6_0_33, w_stg_6_1_33, w_stg_6_2_33);
	assign w_stg_7_2_33 = w_stg_6_3_33;
	full_adder_md fa881( w_stg_7_1_34, w_stg_7_0_35, w_stg_6_0_34, w_stg_6_1_34, w_stg_6_2_34);
	assign w_stg_7_2_34 = w_stg_6_3_34;
	full_adder_md fa882( w_stg_7_1_35, w_stg_7_0_36, w_stg_6_0_35, w_stg_6_1_35, w_stg_6_2_35);
	assign w_stg_7_2_35 = w_stg_6_3_35;
	full_adder_md fa883( w_stg_7_1_36, w_stg_7_0_37, w_stg_6_0_36, w_stg_6_1_36, w_stg_6_2_36);
	assign w_stg_7_2_36 = w_stg_6_3_36;
	full_adder_md fa884( w_stg_7_1_37, w_stg_7_0_38, w_stg_6_0_37, w_stg_6_1_37, w_stg_6_2_37);
	assign w_stg_7_2_37 = w_stg_6_3_37;
	full_adder_md fa885( w_stg_7_1_38, w_stg_7_0_39, w_stg_6_0_38, w_stg_6_1_38, w_stg_6_2_38);
	assign w_stg_7_2_38 = w_stg_6_3_38;
	full_adder_md fa886( w_stg_7_1_39, w_stg_7_0_40, w_stg_6_0_39, w_stg_6_1_39, w_stg_6_2_39);
	full_adder_md fa887( w_stg_7_1_40, w_stg_7_0_41, w_stg_6_0_40, w_stg_6_1_40, w_stg_6_2_40);
	full_adder_md fa888( w_stg_7_1_41, w_stg_7_0_42, w_stg_6_0_41, w_stg_6_1_41, w_stg_6_2_41);
	full_adder_md fa889( w_stg_7_1_42, w_stg_7_0_43, w_stg_6_0_42, w_stg_6_1_42, w_stg_6_2_42);
	full_adder_md fa890( w_stg_7_1_43, w_stg_7_0_44, w_stg_6_0_43, w_stg_6_1_43, w_stg_6_2_43);
	full_adder_md fa891( w_stg_7_1_44, w_stg_7_0_45, w_stg_6_0_44, w_stg_6_1_44, w_stg_6_2_44);
	full_adder_md fa892( w_stg_7_1_45, w_stg_7_0_46, w_stg_6_0_45, w_stg_6_1_45, w_stg_6_2_45);
	full_adder_md fa893( w_stg_7_1_46, w_stg_7_0_47, w_stg_6_0_46, w_stg_6_1_46, w_stg_6_2_46);
	half_adder ha176( w_stg_7_1_47, w_stg_7_0_48, w_stg_6_0_47, w_stg_6_1_47);
	half_adder ha177( w_stg_7_1_48, w_stg_7_0_49, w_stg_6_0_48, w_stg_6_1_48);
	half_adder ha178( w_stg_7_1_49, w_stg_7_0_50, w_stg_6_0_49, w_stg_6_1_49);
	half_adder ha179( w_stg_7_1_50, w_stg_7_0_51, w_stg_6_0_50, w_stg_6_1_50);
	half_adder ha180( w_stg_7_1_51, w_stg_7_0_52, w_stg_6_0_51, w_stg_6_1_51);
	half_adder ha181( w_stg_7_1_52, w_stg_7_0_53, w_stg_6_0_52, w_stg_6_1_52);
	half_adder ha182( w_stg_7_1_53, w_stg_7_0_54, w_stg_6_0_53, w_stg_6_1_53);
	half_adder ha183( w_stg_7_1_54, w_stg_7_0_55, w_stg_6_0_54, w_stg_6_1_54);
	half_adder ha184( w_stg_7_1_55, w_stg_7_0_56, w_stg_6_0_55, w_stg_6_1_55);
	half_adder ha185( w_stg_7_1_56, w_stg_7_0_57, w_stg_6_0_56, w_stg_6_1_56);
	half_adder ha186( w_stg_7_1_57, w_stg_7_0_58, w_stg_6_0_57, w_stg_6_1_57);
	half_adder ha187( w_stg_7_1_58, w_stg_7_0_59, w_stg_6_0_58, w_stg_6_1_58);
	half_adder ha188( w_stg_7_1_59, w_stg_7_0_60, w_stg_6_0_59, w_stg_6_1_59);
	half_adder ha189( w_stg_7_1_60, w_stg_7_0_61, w_stg_6_0_60, w_stg_6_1_60);
	half_adder ha190( w_stg_7_1_61, w_stg_7_0_62, w_stg_6_0_61, w_stg_6_1_61);
	half_adder ha191( w_stg_7_1_62, w_stg_7_0_63, w_stg_6_0_62, w_stg_6_1_62);
	half_adder ha192( w_stg_7_1_63, w_stg_7_0_64, w_stg_6_0_63, w_stg_6_1_63);
	half_adder ha193( w_stg_7_1_64, w_stg_7_0_65, w_stg_6_0_64, w_stg_6_1_64);
	assign w_stg_7_1_65 = w_stg_6_0_65;
	assign w_stg_8_0_0 = w_stg_7_0_0;
	assign w_stg_8_0_1 = w_stg_7_0_1;
	assign w_stg_8_0_2 = w_stg_7_0_2;
	assign w_stg_8_0_3 = w_stg_7_0_3;
	assign w_stg_8_0_4 = w_stg_7_0_4;
	assign w_stg_8_0_5 = w_stg_7_0_5;
	assign w_stg_8_0_6 = w_stg_7_0_6;
	assign w_stg_8_0_7 = w_stg_7_0_7;
	half_adder ha194( w_stg_8_0_8, w_stg_8_0_9, w_stg_7_0_8, w_stg_7_1_8);
	half_adder ha195( w_stg_8_1_9, w_stg_8_0_10, w_stg_7_0_9, w_stg_7_1_9);
	half_adder ha196( w_stg_8_1_10, w_stg_8_0_11, w_stg_7_0_10, w_stg_7_1_10);
	half_adder ha197( w_stg_8_1_11, w_stg_8_0_12, w_stg_7_0_11, w_stg_7_1_11);
	half_adder ha198( w_stg_8_1_12, w_stg_8_0_13, w_stg_7_0_12, w_stg_7_1_12);
	half_adder ha199( w_stg_8_1_13, w_stg_8_0_14, w_stg_7_0_13, w_stg_7_1_13);
	half_adder ha200( w_stg_8_1_14, w_stg_8_0_15, w_stg_7_0_14, w_stg_7_1_14);
	half_adder ha201( w_stg_8_1_15, w_stg_8_0_16, w_stg_7_0_15, w_stg_7_1_15);
	half_adder ha202( w_stg_8_1_16, w_stg_8_0_17, w_stg_7_0_16, w_stg_7_1_16);
	half_adder ha203( w_stg_8_1_17, w_stg_8_0_18, w_stg_7_0_17, w_stg_7_1_17);
	half_adder ha204( w_stg_8_1_18, w_stg_8_0_19, w_stg_7_0_18, w_stg_7_1_18);
	half_adder ha205( w_stg_8_1_19, w_stg_8_0_20, w_stg_7_0_19, w_stg_7_1_19);
	half_adder ha206( w_stg_8_1_20, w_stg_8_0_21, w_stg_7_0_20, w_stg_7_1_20);
	half_adder ha207( w_stg_8_1_21, w_stg_8_0_22, w_stg_7_0_21, w_stg_7_1_21);
	half_adder ha208( w_stg_8_1_22, w_stg_8_0_23, w_stg_7_0_22, w_stg_7_1_22);
	half_adder ha209( w_stg_8_1_23, w_stg_8_0_24, w_stg_7_0_23, w_stg_7_1_23);
	half_adder ha210( w_stg_8_1_24, w_stg_8_0_25, w_stg_7_0_24, w_stg_7_1_24);
	half_adder ha211( w_stg_8_1_25, w_stg_8_0_26, w_stg_7_0_25, w_stg_7_1_25);
	half_adder ha212( w_stg_8_1_26, w_stg_8_0_27, w_stg_7_0_26, w_stg_7_1_26);
	half_adder ha213( w_stg_8_1_27, w_stg_8_0_28, w_stg_7_0_27, w_stg_7_1_27);
	half_adder ha214( w_stg_8_1_28, w_stg_8_0_29, w_stg_7_0_28, w_stg_7_1_28);
	half_adder ha215( w_stg_8_1_29, w_stg_8_0_30, w_stg_7_0_29, w_stg_7_1_29);
	half_adder ha216( w_stg_8_1_30, w_stg_8_0_31, w_stg_7_0_30, w_stg_7_1_30);
	half_adder ha217( w_stg_8_1_31, w_stg_8_0_32, w_stg_7_0_31, w_stg_7_1_31);
	full_adder_md fa894( w_stg_8_1_32, w_stg_8_0_33, w_stg_7_0_32, w_stg_7_1_32, w_stg_7_2_32);
	full_adder_md fa895( w_stg_8_1_33, w_stg_8_0_34, w_stg_7_0_33, w_stg_7_1_33, w_stg_7_2_33);
	full_adder_md fa896( w_stg_8_1_34, w_stg_8_0_35, w_stg_7_0_34, w_stg_7_1_34, w_stg_7_2_34);
	full_adder_md fa897( w_stg_8_1_35, w_stg_8_0_36, w_stg_7_0_35, w_stg_7_1_35, w_stg_7_2_35);
	full_adder_md fa898( w_stg_8_1_36, w_stg_8_0_37, w_stg_7_0_36, w_stg_7_1_36, w_stg_7_2_36);
	full_adder_md fa899( w_stg_8_1_37, w_stg_8_0_38, w_stg_7_0_37, w_stg_7_1_37, w_stg_7_2_37);
	full_adder_md fa900( w_stg_8_1_38, w_stg_8_0_39, w_stg_7_0_38, w_stg_7_1_38, w_stg_7_2_38);
	half_adder ha218( w_stg_8_1_39, w_stg_8_0_40, w_stg_7_0_39, w_stg_7_1_39);
	half_adder ha219( w_stg_8_1_40, w_stg_8_0_41, w_stg_7_0_40, w_stg_7_1_40);
	half_adder ha220( w_stg_8_1_41, w_stg_8_0_42, w_stg_7_0_41, w_stg_7_1_41);
	half_adder ha221( w_stg_8_1_42, w_stg_8_0_43, w_stg_7_0_42, w_stg_7_1_42);
	half_adder ha222( w_stg_8_1_43, w_stg_8_0_44, w_stg_7_0_43, w_stg_7_1_43);
	half_adder ha223( w_stg_8_1_44, w_stg_8_0_45, w_stg_7_0_44, w_stg_7_1_44);
	half_adder ha224( w_stg_8_1_45, w_stg_8_0_46, w_stg_7_0_45, w_stg_7_1_45);
	half_adder ha225( w_stg_8_1_46, w_stg_8_0_47, w_stg_7_0_46, w_stg_7_1_46);
	half_adder ha226( w_stg_8_1_47, w_stg_8_0_48, w_stg_7_0_47, w_stg_7_1_47);
	half_adder ha227( w_stg_8_1_48, w_stg_8_0_49, w_stg_7_0_48, w_stg_7_1_48);
	half_adder ha228( w_stg_8_1_49, w_stg_8_0_50, w_stg_7_0_49, w_stg_7_1_49);
	half_adder ha229( w_stg_8_1_50, w_stg_8_0_51, w_stg_7_0_50, w_stg_7_1_50);
	half_adder ha230( w_stg_8_1_51, w_stg_8_0_52, w_stg_7_0_51, w_stg_7_1_51);
	half_adder ha231( w_stg_8_1_52, w_stg_8_0_53, w_stg_7_0_52, w_stg_7_1_52);
	half_adder ha232( w_stg_8_1_53, w_stg_8_0_54, w_stg_7_0_53, w_stg_7_1_53);
	half_adder ha233( w_stg_8_1_54, w_stg_8_0_55, w_stg_7_0_54, w_stg_7_1_54);
	half_adder ha234( w_stg_8_1_55, w_stg_8_0_56, w_stg_7_0_55, w_stg_7_1_55);
	half_adder ha235( w_stg_8_1_56, w_stg_8_0_57, w_stg_7_0_56, w_stg_7_1_56);
	half_adder ha236( w_stg_8_1_57, w_stg_8_0_58, w_stg_7_0_57, w_stg_7_1_57);
	half_adder ha237( w_stg_8_1_58, w_stg_8_0_59, w_stg_7_0_58, w_stg_7_1_58);
	half_adder ha238( w_stg_8_1_59, w_stg_8_0_60, w_stg_7_0_59, w_stg_7_1_59);
	half_adder ha239( w_stg_8_1_60, w_stg_8_0_61, w_stg_7_0_60, w_stg_7_1_60);
	half_adder ha240( w_stg_8_1_61, w_stg_8_0_62, w_stg_7_0_61, w_stg_7_1_61);
	half_adder ha241( w_stg_8_1_62, w_stg_8_0_63, w_stg_7_0_62, w_stg_7_1_62);
	half_adder ha242( w_stg_8_1_63, w_stg_8_0_64, w_stg_7_0_63, w_stg_7_1_63);
	half_adder ha243( w_stg_8_1_64, w_stg_8_0_65, w_stg_7_0_64, w_stg_7_1_64);
	half_adder ha244( w_stg_8_1_65, w_stg_8_0_66, w_stg_7_0_65, w_stg_7_1_65);

	wire [63:0] x, y;

	assign y[0] = 1'b0;
	assign x[0] = w_stg_8_0_0;
	assign y[1] = 1'b0;
	assign x[1] = w_stg_8_0_1;
	assign y[2] = 1'b0;
	assign x[2] = w_stg_8_0_2;
	assign y[3] = 1'b0;
	assign x[3] = w_stg_8_0_3;
	assign y[4] = 1'b0;
	assign x[4] = w_stg_8_0_4;
	assign y[5] = 1'b0;
	assign x[5] = w_stg_8_0_5;
	assign y[6] = 1'b0;
	assign x[6] = w_stg_8_0_6;
	assign y[7] = 1'b0;
	assign x[7] = w_stg_8_0_7;
	assign y[8] = 1'b0;
	assign x[8] = w_stg_8_0_8;
	assign y[9] = w_stg_8_1_9;
	assign x[9] = w_stg_8_0_9;
	assign y[10] = w_stg_8_1_10;
	assign x[10] = w_stg_8_0_10;
	assign y[11] = w_stg_8_1_11;
	assign x[11] = w_stg_8_0_11;
	assign y[12] = w_stg_8_1_12;
	assign x[12] = w_stg_8_0_12;
	assign y[13] = w_stg_8_1_13;
	assign x[13] = w_stg_8_0_13;
	assign y[14] = w_stg_8_1_14;
	assign x[14] = w_stg_8_0_14;
	assign y[15] = w_stg_8_1_15;
	assign x[15] = w_stg_8_0_15;
	assign y[16] = w_stg_8_1_16;
	assign x[16] = w_stg_8_0_16;
	assign y[17] = w_stg_8_1_17;
	assign x[17] = w_stg_8_0_17;
	assign y[18] = w_stg_8_1_18;
	assign x[18] = w_stg_8_0_18;
	assign y[19] = w_stg_8_1_19;
	assign x[19] = w_stg_8_0_19;
	assign y[20] = w_stg_8_1_20;
	assign x[20] = w_stg_8_0_20;
	assign y[21] = w_stg_8_1_21;
	assign x[21] = w_stg_8_0_21;
	assign y[22] = w_stg_8_1_22;
	assign x[22] = w_stg_8_0_22;
	assign y[23] = w_stg_8_1_23;
	assign x[23] = w_stg_8_0_23;
	assign y[24] = w_stg_8_1_24;
	assign x[24] = w_stg_8_0_24;
	assign y[25] = w_stg_8_1_25;
	assign x[25] = w_stg_8_0_25;
	assign y[26] = w_stg_8_1_26;
	assign x[26] = w_stg_8_0_26;
	assign y[27] = w_stg_8_1_27;
	assign x[27] = w_stg_8_0_27;
	assign y[28] = w_stg_8_1_28;
	assign x[28] = w_stg_8_0_28;
	assign y[29] = w_stg_8_1_29;
	assign x[29] = w_stg_8_0_29;
	assign y[30] = w_stg_8_1_30;
	assign x[30] = w_stg_8_0_30;
	assign y[31] = w_stg_8_1_31;
	assign x[31] = w_stg_8_0_31;
	assign y[32] = w_stg_8_1_32;
	assign x[32] = w_stg_8_0_32;
	assign y[33] = w_stg_8_1_33;
	assign x[33] = w_stg_8_0_33;
	assign y[34] = w_stg_8_1_34;
	assign x[34] = w_stg_8_0_34;
	assign y[35] = w_stg_8_1_35;
	assign x[35] = w_stg_8_0_35;
	assign y[36] = w_stg_8_1_36;
	assign x[36] = w_stg_8_0_36;
	assign y[37] = w_stg_8_1_37;
	assign x[37] = w_stg_8_0_37;
	assign y[38] = w_stg_8_1_38;
	assign x[38] = w_stg_8_0_38;
	assign y[39] = w_stg_8_1_39;
	assign x[39] = w_stg_8_0_39;
	assign y[40] = w_stg_8_1_40;
	assign x[40] = w_stg_8_0_40;
	assign y[41] = w_stg_8_1_41;
	assign x[41] = w_stg_8_0_41;
	assign y[42] = w_stg_8_1_42;
	assign x[42] = w_stg_8_0_42;
	assign y[43] = w_stg_8_1_43;
	assign x[43] = w_stg_8_0_43;
	assign y[44] = w_stg_8_1_44;
	assign x[44] = w_stg_8_0_44;
	assign y[45] = w_stg_8_1_45;
	assign x[45] = w_stg_8_0_45;
	assign y[46] = w_stg_8_1_46;
	assign x[46] = w_stg_8_0_46;
	assign y[47] = w_stg_8_1_47;
	assign x[47] = w_stg_8_0_47;
	assign y[48] = w_stg_8_1_48;
	assign x[48] = w_stg_8_0_48;
	assign y[49] = w_stg_8_1_49;
	assign x[49] = w_stg_8_0_49;
	assign y[50] = w_stg_8_1_50;
	assign x[50] = w_stg_8_0_50;
	assign y[51] = w_stg_8_1_51;
	assign x[51] = w_stg_8_0_51;
	assign y[52] = w_stg_8_1_52;
	assign x[52] = w_stg_8_0_52;
	assign y[53] = w_stg_8_1_53;
	assign x[53] = w_stg_8_0_53;
	assign y[54] = w_stg_8_1_54;
	assign x[54] = w_stg_8_0_54;
	assign y[55] = w_stg_8_1_55;
	assign x[55] = w_stg_8_0_55;
	assign y[56] = w_stg_8_1_56;
	assign x[56] = w_stg_8_0_56;
	assign y[57] = w_stg_8_1_57;
	assign x[57] = w_stg_8_0_57;
	assign y[58] = w_stg_8_1_58;
	assign x[58] = w_stg_8_0_58;
	assign y[59] = w_stg_8_1_59;
	assign x[59] = w_stg_8_0_59;
	assign y[60] = w_stg_8_1_60;
	assign x[60] = w_stg_8_0_60;
	assign y[61] = w_stg_8_1_61;
	assign x[61] = w_stg_8_0_61;
	assign y[62] = w_stg_8_1_62;
	assign x[62] = w_stg_8_0_62;
	assign y[63] = w_stg_8_1_63;
	assign x[63] = w_stg_8_0_63;



	wire [63:0] long_sum;
	wire cout_s1, cout_s2;
	cselect_adder_32 cs1(x[31:0], y[31:0], 1'b0, cout_s1, long_sum[31:0]);
	cselect_adder_32 cs2(x[63:32], y[63:32], cout_s1, cout_s2, long_sum[63:32]);

	assign data_result = long_sum[31:0];
endmodule
