module x_mult(a, b, result, data_exception);
input [31:0] a, b;
output [31:0] result;
output data_exception;
wire [63:0] out1, out2;

wire wand31_0, wand30_0, wand29_0, wand28_0, wand27_0, wand26_0, wand25_0, wand24_0, wand23_0, wand22_0, wand21_0, wand20_0, wand19_0, wand18_0, wand17_0, wand16_0, wand15_0, wand14_0, wand13_0, wand12_0, wand11_0, wand10_0, wand9_0, wand8_0, wand7_0, wand6_0, wand5_0, wand4_0, wand3_0, wand2_0, wand1_0, wand0_0, wand31_1, wand30_1, wand29_1, wand28_1, wand27_1, wand26_1, wand25_1, wand24_1, wand23_1, wand22_1, wand21_1, wand20_1, wand19_1, wand18_1, wand17_1, wand16_1, wand15_1, wand14_1, wand13_1, wand12_1, wand11_1, wand10_1, wand9_1, wand8_1, wand7_1, wand6_1, wand5_1, wand4_1, wand3_1, wand2_1, wand1_1, wand0_1, wand31_2, wand30_2, wand29_2, wand28_2, wand27_2, wand26_2, wand25_2, wand24_2, wand23_2, wand22_2, wand21_2, wand20_2, wand19_2, wand18_2, wand17_2, wand16_2, wand15_2, wand14_2, wand13_2, wand12_2, wand11_2, wand10_2, wand9_2, wand8_2, wand7_2, wand6_2, wand5_2, wand4_2, wand3_2, wand2_2, wand1_2, wand0_2, wand31_3, wand30_3, wand29_3, wand28_3, wand27_3, wand26_3, wand25_3, wand24_3, wand23_3, wand22_3, wand21_3, wand20_3, wand19_3, wand18_3, wand17_3, wand16_3, wand15_3, wand14_3, wand13_3, wand12_3, wand11_3, wand10_3, wand9_3, wand8_3, wand7_3, wand6_3, wand5_3, wand4_3, wand3_3, wand2_3, wand1_3, wand0_3, wand31_4, wand30_4, wand29_4, wand28_4, wand27_4, wand26_4, wand25_4, wand24_4, wand23_4, wand22_4, wand21_4, wand20_4, wand19_4, wand18_4, wand17_4, wand16_4, wand15_4, wand14_4, wand13_4, wand12_4, wand11_4, wand10_4, wand9_4, wand8_4, wand7_4, wand6_4, wand5_4, wand4_4, wand3_4, wand2_4, wand1_4, wand0_4, wand31_5, wand30_5, wand29_5, wand28_5, wand27_5, wand26_5, wand25_5, wand24_5, wand23_5, wand22_5, wand21_5, wand20_5, wand19_5, wand18_5, wand17_5, wand16_5, wand15_5, wand14_5, wand13_5, wand12_5, wand11_5, wand10_5, wand9_5, wand8_5, wand7_5, wand6_5, wand5_5, wand4_5, wand3_5, wand2_5, wand1_5, wand0_5, wand31_6, wand30_6, wand29_6, wand28_6, wand27_6, wand26_6, wand25_6, wand24_6, wand23_6, wand22_6, wand21_6, wand20_6, wand19_6, wand18_6, wand17_6, wand16_6, wand15_6, wand14_6, wand13_6, wand12_6, wand11_6, wand10_6, wand9_6, wand8_6, wand7_6, wand6_6, wand5_6, wand4_6, wand3_6, wand2_6, wand1_6, wand0_6, wand31_7, wand30_7, wand29_7, wand28_7, wand27_7, wand26_7, wand25_7, wand24_7, wand23_7, wand22_7, wand21_7, wand20_7, wand19_7, wand18_7, wand17_7, wand16_7, wand15_7, wand14_7, wand13_7, wand12_7, wand11_7, wand10_7, wand9_7, wand8_7, wand7_7, wand6_7, wand5_7, wand4_7, wand3_7, wand2_7, wand1_7, wand0_7, wand31_8, wand30_8, wand29_8, wand28_8, wand27_8, wand26_8, wand25_8, wand24_8, wand23_8, wand22_8, wand21_8, wand20_8, wand19_8, wand18_8, wand17_8, wand16_8, wand15_8, wand14_8, wand13_8, wand12_8, wand11_8, wand10_8, wand9_8, wand8_8, wand7_8, wand6_8, wand5_8, wand4_8, wand3_8, wand2_8, wand1_8, wand0_8, wand31_9, wand30_9, wand29_9, wand28_9, wand27_9, wand26_9, wand25_9, wand24_9, wand23_9, wand22_9, wand21_9, wand20_9, wand19_9, wand18_9, wand17_9, wand16_9, wand15_9, wand14_9, wand13_9, wand12_9, wand11_9, wand10_9, wand9_9, wand8_9, wand7_9, wand6_9, wand5_9, wand4_9, wand3_9, wand2_9, wand1_9, wand0_9, wand31_10, wand30_10, wand29_10, wand28_10, wand27_10, wand26_10, wand25_10, wand24_10, wand23_10, wand22_10, wand21_10, wand20_10, wand19_10, wand18_10, wand17_10, wand16_10, wand15_10, wand14_10, wand13_10, wand12_10, wand11_10, wand10_10, wand9_10, wand8_10, wand7_10, wand6_10, wand5_10, wand4_10, wand3_10, wand2_10, wand1_10, wand0_10, wand31_11, wand30_11, wand29_11, wand28_11, wand27_11, wand26_11, wand25_11, wand24_11, wand23_11, wand22_11, wand21_11, wand20_11, wand19_11, wand18_11, wand17_11, wand16_11, wand15_11, wand14_11, wand13_11, wand12_11, wand11_11, wand10_11, wand9_11, wand8_11, wand7_11, wand6_11, wand5_11, wand4_11, wand3_11, wand2_11, wand1_11, wand0_11, wand31_12, wand30_12, wand29_12, wand28_12, wand27_12, wand26_12, wand25_12, wand24_12, wand23_12, wand22_12, wand21_12, wand20_12, wand19_12, wand18_12, wand17_12, wand16_12, wand15_12, wand14_12, wand13_12, wand12_12, wand11_12, wand10_12, wand9_12, wand8_12, wand7_12, wand6_12, wand5_12, wand4_12, wand3_12, wand2_12, wand1_12, wand0_12, wand31_13, wand30_13, wand29_13, wand28_13, wand27_13, wand26_13, wand25_13, wand24_13, wand23_13, wand22_13, wand21_13, wand20_13, wand19_13, wand18_13, wand17_13, wand16_13, wand15_13, wand14_13, wand13_13, wand12_13, wand11_13, wand10_13, wand9_13, wand8_13, wand7_13, wand6_13, wand5_13, wand4_13, wand3_13, wand2_13, wand1_13, wand0_13, wand31_14, wand30_14, wand29_14, wand28_14, wand27_14, wand26_14, wand25_14, wand24_14, wand23_14, wand22_14, wand21_14, wand20_14, wand19_14, wand18_14, wand17_14, wand16_14, wand15_14, wand14_14, wand13_14, wand12_14, wand11_14, wand10_14, wand9_14, wand8_14, wand7_14, wand6_14, wand5_14, wand4_14, wand3_14, wand2_14, wand1_14, wand0_14, wand31_15, wand30_15, wand29_15, wand28_15, wand27_15, wand26_15, wand25_15, wand24_15, wand23_15, wand22_15, wand21_15, wand20_15, wand19_15, wand18_15, wand17_15, wand16_15, wand15_15, wand14_15, wand13_15, wand12_15, wand11_15, wand10_15, wand9_15, wand8_15, wand7_15, wand6_15, wand5_15, wand4_15, wand3_15, wand2_15, wand1_15, wand0_15, wand31_16, wand30_16, wand29_16, wand28_16, wand27_16, wand26_16, wand25_16, wand24_16, wand23_16, wand22_16, wand21_16, wand20_16, wand19_16, wand18_16, wand17_16, wand16_16, wand15_16, wand14_16, wand13_16, wand12_16, wand11_16, wand10_16, wand9_16, wand8_16, wand7_16, wand6_16, wand5_16, wand4_16, wand3_16, wand2_16, wand1_16, wand0_16, wand31_17, wand30_17, wand29_17, wand28_17, wand27_17, wand26_17, wand25_17, wand24_17, wand23_17, wand22_17, wand21_17, wand20_17, wand19_17, wand18_17, wand17_17, wand16_17, wand15_17, wand14_17, wand13_17, wand12_17, wand11_17, wand10_17, wand9_17, wand8_17, wand7_17, wand6_17, wand5_17, wand4_17, wand3_17, wand2_17, wand1_17, wand0_17, wand31_18, wand30_18, wand29_18, wand28_18, wand27_18, wand26_18, wand25_18, wand24_18, wand23_18, wand22_18, wand21_18, wand20_18, wand19_18, wand18_18, wand17_18, wand16_18, wand15_18, wand14_18, wand13_18, wand12_18, wand11_18, wand10_18, wand9_18, wand8_18, wand7_18, wand6_18, wand5_18, wand4_18, wand3_18, wand2_18, wand1_18, wand0_18, wand31_19, wand30_19, wand29_19, wand28_19, wand27_19, wand26_19, wand25_19, wand24_19, wand23_19, wand22_19, wand21_19, wand20_19, wand19_19, wand18_19, wand17_19, wand16_19, wand15_19, wand14_19, wand13_19, wand12_19, wand11_19, wand10_19, wand9_19, wand8_19, wand7_19, wand6_19, wand5_19, wand4_19, wand3_19, wand2_19, wand1_19, wand0_19, wand31_20, wand30_20, wand29_20, wand28_20, wand27_20, wand26_20, wand25_20, wand24_20, wand23_20, wand22_20, wand21_20, wand20_20, wand19_20, wand18_20, wand17_20, wand16_20, wand15_20, wand14_20, wand13_20, wand12_20, wand11_20, wand10_20, wand9_20, wand8_20, wand7_20, wand6_20, wand5_20, wand4_20, wand3_20, wand2_20, wand1_20, wand0_20, wand31_21, wand30_21, wand29_21, wand28_21, wand27_21, wand26_21, wand25_21, wand24_21, wand23_21, wand22_21, wand21_21, wand20_21, wand19_21, wand18_21, wand17_21, wand16_21, wand15_21, wand14_21, wand13_21, wand12_21, wand11_21, wand10_21, wand9_21, wand8_21, wand7_21, wand6_21, wand5_21, wand4_21, wand3_21, wand2_21, wand1_21, wand0_21, wand31_22, wand30_22, wand29_22, wand28_22, wand27_22, wand26_22, wand25_22, wand24_22, wand23_22, wand22_22, wand21_22, wand20_22, wand19_22, wand18_22, wand17_22, wand16_22, wand15_22, wand14_22, wand13_22, wand12_22, wand11_22, wand10_22, wand9_22, wand8_22, wand7_22, wand6_22, wand5_22, wand4_22, wand3_22, wand2_22, wand1_22, wand0_22, wand31_23, wand30_23, wand29_23, wand28_23, wand27_23, wand26_23, wand25_23, wand24_23, wand23_23, wand22_23, wand21_23, wand20_23, wand19_23, wand18_23, wand17_23, wand16_23, wand15_23, wand14_23, wand13_23, wand12_23, wand11_23, wand10_23, wand9_23, wand8_23, wand7_23, wand6_23, wand5_23, wand4_23, wand3_23, wand2_23, wand1_23, wand0_23, wand31_24, wand30_24, wand29_24, wand28_24, wand27_24, wand26_24, wand25_24, wand24_24, wand23_24, wand22_24, wand21_24, wand20_24, wand19_24, wand18_24, wand17_24, wand16_24, wand15_24, wand14_24, wand13_24, wand12_24, wand11_24, wand10_24, wand9_24, wand8_24, wand7_24, wand6_24, wand5_24, wand4_24, wand3_24, wand2_24, wand1_24, wand0_24, wand31_25, wand30_25, wand29_25, wand28_25, wand27_25, wand26_25, wand25_25, wand24_25, wand23_25, wand22_25, wand21_25, wand20_25, wand19_25, wand18_25, wand17_25, wand16_25, wand15_25, wand14_25, wand13_25, wand12_25, wand11_25, wand10_25, wand9_25, wand8_25, wand7_25, wand6_25, wand5_25, wand4_25, wand3_25, wand2_25, wand1_25, wand0_25, wand31_26, wand30_26, wand29_26, wand28_26, wand27_26, wand26_26, wand25_26, wand24_26, wand23_26, wand22_26, wand21_26, wand20_26, wand19_26, wand18_26, wand17_26, wand16_26, wand15_26, wand14_26, wand13_26, wand12_26, wand11_26, wand10_26, wand9_26, wand8_26, wand7_26, wand6_26, wand5_26, wand4_26, wand3_26, wand2_26, wand1_26, wand0_26, wand31_27, wand30_27, wand29_27, wand28_27, wand27_27, wand26_27, wand25_27, wand24_27, wand23_27, wand22_27, wand21_27, wand20_27, wand19_27, wand18_27, wand17_27, wand16_27, wand15_27, wand14_27, wand13_27, wand12_27, wand11_27, wand10_27, wand9_27, wand8_27, wand7_27, wand6_27, wand5_27, wand4_27, wand3_27, wand2_27, wand1_27, wand0_27, wand31_28, wand30_28, wand29_28, wand28_28, wand27_28, wand26_28, wand25_28, wand24_28, wand23_28, wand22_28, wand21_28, wand20_28, wand19_28, wand18_28, wand17_28, wand16_28, wand15_28, wand14_28, wand13_28, wand12_28, wand11_28, wand10_28, wand9_28, wand8_28, wand7_28, wand6_28, wand5_28, wand4_28, wand3_28, wand2_28, wand1_28, wand0_28, wand31_29, wand30_29, wand29_29, wand28_29, wand27_29, wand26_29, wand25_29, wand24_29, wand23_29, wand22_29, wand21_29, wand20_29, wand19_29, wand18_29, wand17_29, wand16_29, wand15_29, wand14_29, wand13_29, wand12_29, wand11_29, wand10_29, wand9_29, wand8_29, wand7_29, wand6_29, wand5_29, wand4_29, wand3_29, wand2_29, wand1_29, wand0_29, wand31_30, wand30_30, wand29_30, wand28_30, wand27_30, wand26_30, wand25_30, wand24_30, wand23_30, wand22_30, wand21_30, wand20_30, wand19_30, wand18_30, wand17_30, wand16_30, wand15_30, wand14_30, wand13_30, wand12_30, wand11_30, wand10_30, wand9_30, wand8_30, wand7_30, wand6_30, wand5_30, wand4_30, wand3_30, wand2_30, wand1_30, wand0_30, wand31_31, wand30_31, wand29_31, wand28_31, wand27_31, wand26_31, wand25_31, wand24_31, wand23_31, wand22_31, wand21_31, wand20_31, wand19_31, wand18_31, wand17_31, wand16_31, wand15_31, wand14_31, wand13_31, wand12_31, wand11_31, wand10_31, wand9_31, wand8_31, wand7_31, wand6_31, wand5_31, wand4_31, wand3_31, wand2_31, wand1_31, wand0_31;
wire ws0b0n0_30, ws0b0n0_31, ws0b0n1_30, ws0b0n0_32, ws0b0n1_31, ws0b0n0_33, ws0b0n1_32, ws0b0n0_34, ws0b0n1_33, ws0b0n0_35, ws0b0n1_34, ws0b0n0_36, ws0b0n1_35, ws0b0n0_37, ws0b0n1_36, ws0b0n0_38, ws0b0n1_37, ws0b0n0_39, ws0b0n1_38, ws0b0n0_40, ws0b0n1_39, ws0b0n0_41, ws0b0n1_40, ws0b0n0_42, ws0b0n1_41, ws0b0n0_43, ws0b0n1_42, ws0b0n0_44, ws0b0n1_43, ws0b0n0_45, ws0b0n1_44, ws0b0n0_46, ws0b0n1_45, ws0b0n0_47, ws0b0n1_46, ws0b0n0_48, ws0b0n1_47, ws0b0n0_49, ws0b0n1_48, ws0b0n0_50, ws0b0n1_49, ws0b0n0_51, ws0b0n1_50, ws0b0n0_52, ws0b0n1_51, ws0b0n0_53, ws0b0n1_52, ws0b0n0_54, ws0b0n1_53, ws0b0n0_55, ws0b0n1_54, ws0b0n0_56, ws0b0n1_55, ws0b0n0_57, ws0b0n1_56, ws0b0n0_58, ws0b0n1_57, ws0b0n0_59, ws0b0n1_58, ws0b0n0_60, ws0b0n1_59, ws0b0n0_61, ws0b0n1_60, ws0b0n0_62, ws0b0n1_61, ws0b0n0_63, ws0b1n0_27, ws0b1n0_28, ws0b1n1_27, ws0b1n0_29, ws0b1n1_28, ws0b1n0_30, ws0b1n1_29, ws0b1n0_31, ws0b1n1_30, ws0b1n0_32, ws0b1n1_31, ws0b1n0_33, ws0b1n1_32, ws0b1n0_34, ws0b1n1_33, ws0b1n0_35, ws0b1n1_34, ws0b1n0_36, ws0b1n1_35, ws0b1n0_37, ws0b1n1_36, ws0b1n0_38, ws0b1n1_37, ws0b1n0_39, ws0b1n1_38, ws0b1n0_40, ws0b1n1_39, ws0b1n0_41, ws0b1n1_40, ws0b1n0_42, ws0b1n1_41, ws0b1n0_43, ws0b1n1_42, ws0b1n0_44, ws0b1n1_43, ws0b1n0_45, ws0b1n1_44, ws0b1n0_46, ws0b1n1_45, ws0b1n0_47, ws0b1n1_46, ws0b1n0_48, ws0b1n1_47, ws0b1n0_49, ws0b1n1_48, ws0b1n0_50, ws0b1n1_49, ws0b1n0_51, ws0b1n1_50, ws0b1n0_52, ws0b1n1_51, ws0b1n0_53, ws0b1n1_52, ws0b1n0_54, ws0b1n1_53, ws0b1n0_55, ws0b1n1_54, ws0b1n0_56, ws0b1n1_55, ws0b1n0_57, ws0b1n1_56, ws0b1n0_58, ws0b1n1_57, ws0b1n0_59, ws0b1n1_58, ws0b1n0_60, ws0b2n0_24, ws0b2n0_25, ws0b2n1_24, ws0b2n0_26, ws0b2n1_25, ws0b2n0_27, ws0b2n1_26, ws0b2n0_28, ws0b2n1_27, ws0b2n0_29, ws0b2n1_28, ws0b2n0_30, ws0b2n1_29, ws0b2n0_31, ws0b2n1_30, ws0b2n0_32, ws0b2n1_31, ws0b2n0_33, ws0b2n1_32, ws0b2n0_34, ws0b2n1_33, ws0b2n0_35, ws0b2n1_34, ws0b2n0_36, ws0b2n1_35, ws0b2n0_37, ws0b2n1_36, ws0b2n0_38, ws0b2n1_37, ws0b2n0_39, ws0b2n1_38, ws0b2n0_40, ws0b2n1_39, ws0b2n0_41, ws0b2n1_40, ws0b2n0_42, ws0b2n1_41, ws0b2n0_43, ws0b2n1_42, ws0b2n0_44, ws0b2n1_43, ws0b2n0_45, ws0b2n1_44, ws0b2n0_46, ws0b2n1_45, ws0b2n0_47, ws0b2n1_46, ws0b2n0_48, ws0b2n1_47, ws0b2n0_49, ws0b2n1_48, ws0b2n0_50, ws0b2n1_49, ws0b2n0_51, ws0b2n1_50, ws0b2n0_52, ws0b2n1_51, ws0b2n0_53, ws0b2n1_52, ws0b2n0_54, ws0b2n1_53, ws0b2n0_55, ws0b2n1_54, ws0b2n0_56, ws0b2n1_55, ws0b2n0_57, ws0b3n0_21, ws0b3n0_22, ws0b3n1_21, ws0b3n0_23, ws0b3n1_22, ws0b3n0_24, ws0b3n1_23, ws0b3n0_25, ws0b3n1_24, ws0b3n0_26, ws0b3n1_25, ws0b3n0_27, ws0b3n1_26, ws0b3n0_28, ws0b3n1_27, ws0b3n0_29, ws0b3n1_28, ws0b3n0_30, ws0b3n1_29, ws0b3n0_31, ws0b3n1_30, ws0b3n0_32, ws0b3n1_31, ws0b3n0_33, ws0b3n1_32, ws0b3n0_34, ws0b3n1_33, ws0b3n0_35, ws0b3n1_34, ws0b3n0_36, ws0b3n1_35, ws0b3n0_37, ws0b3n1_36, ws0b3n0_38, ws0b3n1_37, ws0b3n0_39, ws0b3n1_38, ws0b3n0_40, ws0b3n1_39, ws0b3n0_41, ws0b3n1_40, ws0b3n0_42, ws0b3n1_41, ws0b3n0_43, ws0b3n1_42, ws0b3n0_44, ws0b3n1_43, ws0b3n0_45, ws0b3n1_44, ws0b3n0_46, ws0b3n1_45, ws0b3n0_47, ws0b3n1_46, ws0b3n0_48, ws0b3n1_47, ws0b3n0_49, ws0b3n1_48, ws0b3n0_50, ws0b3n1_49, ws0b3n0_51, ws0b3n1_50, ws0b3n0_52, ws0b3n1_51, ws0b3n0_53, ws0b3n1_52, ws0b3n0_54, ws0b4n0_18, ws0b4n0_19, ws0b4n1_18, ws0b4n0_20, ws0b4n1_19, ws0b4n0_21, ws0b4n1_20, ws0b4n0_22, ws0b4n1_21, ws0b4n0_23, ws0b4n1_22, ws0b4n0_24, ws0b4n1_23, ws0b4n0_25, ws0b4n1_24, ws0b4n0_26, ws0b4n1_25, ws0b4n0_27, ws0b4n1_26, ws0b4n0_28, ws0b4n1_27, ws0b4n0_29, ws0b4n1_28, ws0b4n0_30, ws0b4n1_29, ws0b4n0_31, ws0b4n1_30, ws0b4n0_32, ws0b4n1_31, ws0b4n0_33, ws0b4n1_32, ws0b4n0_34, ws0b4n1_33, ws0b4n0_35, ws0b4n1_34, ws0b4n0_36, ws0b4n1_35, ws0b4n0_37, ws0b4n1_36, ws0b4n0_38, ws0b4n1_37, ws0b4n0_39, ws0b4n1_38, ws0b4n0_40, ws0b4n1_39, ws0b4n0_41, ws0b4n1_40, ws0b4n0_42, ws0b4n1_41, ws0b4n0_43, ws0b4n1_42, ws0b4n0_44, ws0b4n1_43, ws0b4n0_45, ws0b4n1_44, ws0b4n0_46, ws0b4n1_45, ws0b4n0_47, ws0b4n1_46, ws0b4n0_48, ws0b4n1_47, ws0b4n0_49, ws0b4n1_48, ws0b4n0_50, ws0b4n1_49, ws0b4n0_51, ws0b5n0_15, ws0b5n0_16, ws0b5n1_15, ws0b5n0_17, ws0b5n1_16, ws0b5n0_18, ws0b5n1_17, ws0b5n0_19, ws0b5n1_18, ws0b5n0_20, ws0b5n1_19, ws0b5n0_21, ws0b5n1_20, ws0b5n0_22, ws0b5n1_21, ws0b5n0_23, ws0b5n1_22, ws0b5n0_24, ws0b5n1_23, ws0b5n0_25, ws0b5n1_24, ws0b5n0_26, ws0b5n1_25, ws0b5n0_27, ws0b5n1_26, ws0b5n0_28, ws0b5n1_27, ws0b5n0_29, ws0b5n1_28, ws0b5n0_30, ws0b5n1_29, ws0b5n0_31, ws0b5n1_30, ws0b5n0_32, ws0b5n1_31, ws0b5n0_33, ws0b5n1_32, ws0b5n0_34, ws0b5n1_33, ws0b5n0_35, ws0b5n1_34, ws0b5n0_36, ws0b5n1_35, ws0b5n0_37, ws0b5n1_36, ws0b5n0_38, ws0b5n1_37, ws0b5n0_39, ws0b5n1_38, ws0b5n0_40, ws0b5n1_39, ws0b5n0_41, ws0b5n1_40, ws0b5n0_42, ws0b5n1_41, ws0b5n0_43, ws0b5n1_42, ws0b5n0_44, ws0b5n1_43, ws0b5n0_45, ws0b5n1_44, ws0b5n0_46, ws0b5n1_45, ws0b5n0_47, ws0b5n1_46, ws0b5n0_48, ws0b6n0_12, ws0b6n0_13, ws0b6n1_12, ws0b6n0_14, ws0b6n1_13, ws0b6n0_15, ws0b6n1_14, ws0b6n0_16, ws0b6n1_15, ws0b6n0_17, ws0b6n1_16, ws0b6n0_18, ws0b6n1_17, ws0b6n0_19, ws0b6n1_18, ws0b6n0_20, ws0b6n1_19, ws0b6n0_21, ws0b6n1_20, ws0b6n0_22, ws0b6n1_21, ws0b6n0_23, ws0b6n1_22, ws0b6n0_24, ws0b6n1_23, ws0b6n0_25, ws0b6n1_24, ws0b6n0_26, ws0b6n1_25, ws0b6n0_27, ws0b6n1_26, ws0b6n0_28, ws0b6n1_27, ws0b6n0_29, ws0b6n1_28, ws0b6n0_30, ws0b6n1_29, ws0b6n0_31, ws0b6n1_30, ws0b6n0_32, ws0b6n1_31, ws0b6n0_33, ws0b6n1_32, ws0b6n0_34, ws0b6n1_33, ws0b6n0_35, ws0b6n1_34, ws0b6n0_36, ws0b6n1_35, ws0b6n0_37, ws0b6n1_36, ws0b6n0_38, ws0b6n1_37, ws0b6n0_39, ws0b6n1_38, ws0b6n0_40, ws0b6n1_39, ws0b6n0_41, ws0b6n1_40, ws0b6n0_42, ws0b6n1_41, ws0b6n0_43, ws0b6n1_42, ws0b6n0_44, ws0b6n1_43, ws0b6n0_45, ws0b7n0_9, ws0b7n0_10, ws0b7n1_9, ws0b7n0_11, ws0b7n1_10, ws0b7n0_12, ws0b7n1_11, ws0b7n0_13, ws0b7n1_12, ws0b7n0_14, ws0b7n1_13, ws0b7n0_15, ws0b7n1_14, ws0b7n0_16, ws0b7n1_15, ws0b7n0_17, ws0b7n1_16, ws0b7n0_18, ws0b7n1_17, ws0b7n0_19, ws0b7n1_18, ws0b7n0_20, ws0b7n1_19, ws0b7n0_21, ws0b7n1_20, ws0b7n0_22, ws0b7n1_21, ws0b7n0_23, ws0b7n1_22, ws0b7n0_24, ws0b7n1_23, ws0b7n0_25, ws0b7n1_24, ws0b7n0_26, ws0b7n1_25, ws0b7n0_27, ws0b7n1_26, ws0b7n0_28, ws0b7n1_27, ws0b7n0_29, ws0b7n1_28, ws0b7n0_30, ws0b7n1_29, ws0b7n0_31, ws0b7n1_30, ws0b7n0_32, ws0b7n1_31, ws0b7n0_33, ws0b7n1_32, ws0b7n0_34, ws0b7n1_33, ws0b7n0_35, ws0b7n1_34, ws0b7n0_36, ws0b7n1_35, ws0b7n0_37, ws0b7n1_36, ws0b7n0_38, ws0b7n1_37, ws0b7n0_39, ws0b7n1_38, ws0b7n0_40, ws0b7n1_39, ws0b7n0_41, ws0b7n1_40, ws0b7n0_42, ws0b8n0_6, ws0b8n0_7, ws0b8n1_6, ws0b8n0_8, ws0b8n1_7, ws0b8n0_9, ws0b8n1_8, ws0b8n0_10, ws0b8n1_9, ws0b8n0_11, ws0b8n1_10, ws0b8n0_12, ws0b8n1_11, ws0b8n0_13, ws0b8n1_12, ws0b8n0_14, ws0b8n1_13, ws0b8n0_15, ws0b8n1_14, ws0b8n0_16, ws0b8n1_15, ws0b8n0_17, ws0b8n1_16, ws0b8n0_18, ws0b8n1_17, ws0b8n0_19, ws0b8n1_18, ws0b8n0_20, ws0b8n1_19, ws0b8n0_21, ws0b8n1_20, ws0b8n0_22, ws0b8n1_21, ws0b8n0_23, ws0b8n1_22, ws0b8n0_24, ws0b8n1_23, ws0b8n0_25, ws0b8n1_24, ws0b8n0_26, ws0b8n1_25, ws0b8n0_27, ws0b8n1_26, ws0b8n0_28, ws0b8n1_27, ws0b8n0_29, ws0b8n1_28, ws0b8n0_30, ws0b8n1_29, ws0b8n0_31, ws0b8n1_30, ws0b8n0_32, ws0b8n1_31, ws0b8n0_33, ws0b8n1_32, ws0b8n0_34, ws0b8n1_33, ws0b8n0_35, ws0b8n1_34, ws0b8n0_36, ws0b8n1_35, ws0b8n0_37, ws0b8n1_36, ws0b8n0_38, ws0b8n1_37, ws0b8n0_39, ws0b9n0_3, ws0b9n0_4, ws0b9n1_3, ws0b9n0_5, ws0b9n1_4, ws0b9n0_6, ws0b9n1_5, ws0b9n0_7, ws0b9n1_6, ws0b9n0_8, ws0b9n1_7, ws0b9n0_9, ws0b9n1_8, ws0b9n0_10, ws0b9n1_9, ws0b9n0_11, ws0b9n1_10, ws0b9n0_12, ws0b9n1_11, ws0b9n0_13, ws0b9n1_12, ws0b9n0_14, ws0b9n1_13, ws0b9n0_15, ws0b9n1_14, ws0b9n0_16, ws0b9n1_15, ws0b9n0_17, ws0b9n1_16, ws0b9n0_18, ws0b9n1_17, ws0b9n0_19, ws0b9n1_18, ws0b9n0_20, ws0b9n1_19, ws0b9n0_21, ws0b9n1_20, ws0b9n0_22, ws0b9n1_21, ws0b9n0_23, ws0b9n1_22, ws0b9n0_24, ws0b9n1_23, ws0b9n0_25, ws0b9n1_24, ws0b9n0_26, ws0b9n1_25, ws0b9n0_27, ws0b9n1_26, ws0b9n0_28, ws0b9n1_27, ws0b9n0_29, ws0b9n1_28, ws0b9n0_30, ws0b9n1_29, ws0b9n0_31, ws0b9n1_30, ws0b9n0_32, ws0b9n1_31, ws0b9n0_33, ws0b9n1_32, ws0b9n0_34, ws0b9n1_33, ws0b9n0_35, ws0b9n1_34, ws0b9n0_36;
wire ws1b0n0_27, ws1b0n0_28, ws1b0n0_29, ws1b0n0_30, ws1b0n1_29, ws1b0n0_31, ws1b0n1_30, ws1b0n0_32, ws1b0n1_31, ws1b0n0_33, ws1b0n1_32, ws1b0n0_34, ws1b0n1_33, ws1b0n0_35, ws1b0n1_34, ws1b0n0_36, ws1b0n1_35, ws1b0n0_37, ws1b0n1_36, ws1b0n0_38, ws1b0n1_37, ws1b0n0_39, ws1b0n1_38, ws1b0n0_40, ws1b0n1_39, ws1b0n0_41, ws1b0n1_40, ws1b0n0_42, ws1b0n1_41, ws1b0n0_43, ws1b0n1_42, ws1b0n0_44, ws1b0n1_43, ws1b0n0_45, ws1b0n1_44, ws1b0n0_46, ws1b0n1_45, ws1b0n0_47, ws1b0n1_46, ws1b0n0_48, ws1b0n1_47, ws1b0n0_49, ws1b0n1_48, ws1b0n0_50, ws1b0n1_49, ws1b0n0_51, ws1b0n1_50, ws1b0n0_52, ws1b0n1_51, ws1b0n0_53, ws1b0n1_52, ws1b0n0_54, ws1b0n1_53, ws1b0n0_55, ws1b0n1_54, ws1b0n0_56, ws1b0n1_55, ws1b0n0_57, ws1b0n1_56, ws1b0n0_58, ws1b0n1_57, ws1b0n0_59, ws1b0n1_58, ws1b0n0_60, ws1b0n1_59, ws1b0n0_61, ws1b0n1_60, ws1b0n0_62, ws1b0n0_63, ws1b1n0_24, ws1b1n1_23, ws1b1n0_25, ws1b1n1_24, ws1b1n0_26, ws1b1n1_25, ws1b1n0_27, ws1b1n1_26, ws1b1n0_28, ws1b1n1_27, ws1b1n0_29, ws1b1n1_28, ws1b1n0_30, ws1b1n1_29, ws1b1n0_31, ws1b1n1_30, ws1b1n0_32, ws1b1n1_31, ws1b1n0_33, ws1b1n1_32, ws1b1n0_34, ws1b1n1_33, ws1b1n0_35, ws1b1n1_34, ws1b1n0_36, ws1b1n1_35, ws1b1n0_37, ws1b1n1_36, ws1b1n0_38, ws1b1n1_37, ws1b1n0_39, ws1b1n1_38, ws1b1n0_40, ws1b1n1_39, ws1b1n0_41, ws1b1n1_40, ws1b1n0_42, ws1b1n1_41, ws1b1n0_43, ws1b1n1_42, ws1b1n0_44, ws1b1n1_43, ws1b1n0_45, ws1b1n1_44, ws1b1n0_46, ws1b1n1_45, ws1b1n0_47, ws1b1n1_46, ws1b1n0_48, ws1b1n1_47, ws1b1n0_49, ws1b1n1_48, ws1b1n0_50, ws1b1n1_49, ws1b1n0_51, ws1b1n1_50, ws1b1n0_52, ws1b1n1_51, ws1b1n0_53, ws1b1n1_52, ws1b1n0_54, ws1b1n1_53, ws1b1n0_55, ws1b1n1_54, ws1b1n0_56, ws1b1n1_55, ws1b1n0_57, ws1b1n1_56, ws1b1n0_58, ws1b2n0_18, ws1b2n0_19, ws1b2n0_20, ws1b2n0_21, ws1b2n1_20, ws1b2n0_22, ws1b2n1_21, ws1b2n0_23, ws1b2n1_22, ws1b2n0_24, ws1b2n1_23, ws1b2n0_25, ws1b2n1_24, ws1b2n0_26, ws1b2n1_25, ws1b2n0_27, ws1b2n1_26, ws1b2n0_28, ws1b2n1_27, ws1b2n0_29, ws1b2n1_28, ws1b2n0_30, ws1b2n1_29, ws1b2n0_31, ws1b2n1_30, ws1b2n0_32, ws1b2n1_31, ws1b2n0_33, ws1b2n1_32, ws1b2n0_34, ws1b2n1_33, ws1b2n0_35, ws1b2n1_34, ws1b2n0_36, ws1b2n1_35, ws1b2n0_37, ws1b2n1_36, ws1b2n0_38, ws1b2n1_37, ws1b2n0_39, ws1b2n1_38, ws1b2n0_40, ws1b2n1_39, ws1b2n0_41, ws1b2n1_40, ws1b2n0_42, ws1b2n1_41, ws1b2n0_43, ws1b2n1_42, ws1b2n0_44, ws1b2n1_43, ws1b2n0_45, ws1b2n1_44, ws1b2n0_46, ws1b2n1_45, ws1b2n0_47, ws1b2n1_46, ws1b2n0_48, ws1b2n1_47, ws1b2n0_49, ws1b2n1_48, ws1b2n0_50, ws1b2n1_49, ws1b2n0_51, ws1b2n1_50, ws1b2n0_52, ws1b2n1_51, ws1b2n0_53, ws1b2n0_54, ws1b3n0_15, ws1b3n1_14, ws1b3n0_16, ws1b3n1_15, ws1b3n0_17, ws1b3n1_16, ws1b3n0_18, ws1b3n1_17, ws1b3n0_19, ws1b3n1_18, ws1b3n0_20, ws1b3n1_19, ws1b3n0_21, ws1b3n1_20, ws1b3n0_22, ws1b3n1_21, ws1b3n0_23, ws1b3n1_22, ws1b3n0_24, ws1b3n1_23, ws1b3n0_25, ws1b3n1_24, ws1b3n0_26, ws1b3n1_25, ws1b3n0_27, ws1b3n1_26, ws1b3n0_28, ws1b3n1_27, ws1b3n0_29, ws1b3n1_28, ws1b3n0_30, ws1b3n1_29, ws1b3n0_31, ws1b3n1_30, ws1b3n0_32, ws1b3n1_31, ws1b3n0_33, ws1b3n1_32, ws1b3n0_34, ws1b3n1_33, ws1b3n0_35, ws1b3n1_34, ws1b3n0_36, ws1b3n1_35, ws1b3n0_37, ws1b3n1_36, ws1b3n0_38, ws1b3n1_37, ws1b3n0_39, ws1b3n1_38, ws1b3n0_40, ws1b3n1_39, ws1b3n0_41, ws1b3n1_40, ws1b3n0_42, ws1b3n1_41, ws1b3n0_43, ws1b3n1_42, ws1b3n0_44, ws1b3n1_43, ws1b3n0_45, ws1b3n1_44, ws1b3n0_46, ws1b3n1_45, ws1b3n0_47, ws1b3n1_46, ws1b3n0_48, ws1b3n1_47, ws1b3n0_49, ws1b4n0_9, ws1b4n0_10, ws1b4n0_11, ws1b4n0_12, ws1b4n1_11, ws1b4n0_13, ws1b4n1_12, ws1b4n0_14, ws1b4n1_13, ws1b4n0_15, ws1b4n1_14, ws1b4n0_16, ws1b4n1_15, ws1b4n0_17, ws1b4n1_16, ws1b4n0_18, ws1b4n1_17, ws1b4n0_19, ws1b4n1_18, ws1b4n0_20, ws1b4n1_19, ws1b4n0_21, ws1b4n1_20, ws1b4n0_22, ws1b4n1_21, ws1b4n0_23, ws1b4n1_22, ws1b4n0_24, ws1b4n1_23, ws1b4n0_25, ws1b4n1_24, ws1b4n0_26, ws1b4n1_25, ws1b4n0_27, ws1b4n1_26, ws1b4n0_28, ws1b4n1_27, ws1b4n0_29, ws1b4n1_28, ws1b4n0_30, ws1b4n1_29, ws1b4n0_31, ws1b4n1_30, ws1b4n0_32, ws1b4n1_31, ws1b4n0_33, ws1b4n1_32, ws1b4n0_34, ws1b4n1_33, ws1b4n0_35, ws1b4n1_34, ws1b4n0_36, ws1b4n1_35, ws1b4n0_37, ws1b4n1_36, ws1b4n0_38, ws1b4n1_37, ws1b4n0_39, ws1b4n1_38, ws1b4n0_40, ws1b4n1_39, ws1b4n0_41, ws1b4n1_40, ws1b4n0_42, ws1b4n1_41, ws1b4n0_43, ws1b4n1_42, ws1b4n0_44, ws1b4n0_45, ws1b5n0_6, ws1b5n1_5, ws1b5n0_7, ws1b5n1_6, ws1b5n0_8, ws1b5n1_7, ws1b5n0_9, ws1b5n1_8, ws1b5n0_10, ws1b5n1_9, ws1b5n0_11, ws1b5n1_10, ws1b5n0_12, ws1b5n1_11, ws1b5n0_13, ws1b5n1_12, ws1b5n0_14, ws1b5n1_13, ws1b5n0_15, ws1b5n1_14, ws1b5n0_16, ws1b5n1_15, ws1b5n0_17, ws1b5n1_16, ws1b5n0_18, ws1b5n1_17, ws1b5n0_19, ws1b5n1_18, ws1b5n0_20, ws1b5n1_19, ws1b5n0_21, ws1b5n1_20, ws1b5n0_22, ws1b5n1_21, ws1b5n0_23, ws1b5n1_22, ws1b5n0_24, ws1b5n1_23, ws1b5n0_25, ws1b5n1_24, ws1b5n0_26, ws1b5n1_25, ws1b5n0_27, ws1b5n1_26, ws1b5n0_28, ws1b5n1_27, ws1b5n0_29, ws1b5n1_28, ws1b5n0_30, ws1b5n1_29, ws1b5n0_31, ws1b5n1_30, ws1b5n0_32, ws1b5n1_31, ws1b5n0_33, ws1b5n1_32, ws1b5n0_34, ws1b5n1_33, ws1b5n0_35, ws1b5n1_34, ws1b5n0_36, ws1b5n1_35, ws1b5n0_37, ws1b5n1_36, ws1b5n0_38, ws1b5n1_37, ws1b5n0_39, ws1b5n1_38, ws1b5n0_40, ws1b6n0_2, ws1b6n0_3, ws1b6n1_2, ws1b6n0_4, ws1b6n1_3, ws1b6n0_5, ws1b6n1_4, ws1b6n0_6, ws1b6n1_5, ws1b6n0_7, ws1b6n1_6, ws1b6n0_8, ws1b6n1_7, ws1b6n0_9, ws1b6n1_8, ws1b6n0_10, ws1b6n1_9, ws1b6n0_11, ws1b6n1_10, ws1b6n0_12, ws1b6n1_11, ws1b6n0_13, ws1b6n1_12, ws1b6n0_14, ws1b6n1_13, ws1b6n0_15, ws1b6n1_14, ws1b6n0_16, ws1b6n1_15, ws1b6n0_17, ws1b6n1_16, ws1b6n0_18, ws1b6n1_17, ws1b6n0_19, ws1b6n1_18, ws1b6n0_20, ws1b6n1_19, ws1b6n0_21, ws1b6n1_20, ws1b6n0_22, ws1b6n1_21, ws1b6n0_23, ws1b6n1_22, ws1b6n0_24, ws1b6n1_23, ws1b6n0_25, ws1b6n1_24, ws1b6n0_26, ws1b6n1_25, ws1b6n0_27, ws1b6n1_26, ws1b6n0_28, ws1b6n1_27, ws1b6n0_29, ws1b6n1_28, ws1b6n0_30, ws1b6n1_29, ws1b6n0_31, ws1b6n1_30, ws1b6n0_32, ws1b6n1_31, ws1b6n0_33, ws1b6n1_32, ws1b6n0_34, ws1b6n1_33, ws1b6n0_35, ws1b6n0_36;
wire ws2b0n0_24, ws2b0n0_25, ws2b0n0_26, ws2b0n0_27, ws2b0n1_26, ws2b0n0_28, ws2b0n1_27, ws2b0n0_29, ws2b0n1_28, ws2b0n0_30, ws2b0n1_29, ws2b0n0_31, ws2b0n1_30, ws2b0n0_32, ws2b0n1_31, ws2b0n0_33, ws2b0n1_32, ws2b0n0_34, ws2b0n1_33, ws2b0n0_35, ws2b0n1_34, ws2b0n0_36, ws2b0n1_35, ws2b0n0_37, ws2b0n1_36, ws2b0n0_38, ws2b0n1_37, ws2b0n0_39, ws2b0n1_38, ws2b0n0_40, ws2b0n1_39, ws2b0n0_41, ws2b0n1_40, ws2b0n0_42, ws2b0n1_41, ws2b0n0_43, ws2b0n1_42, ws2b0n0_44, ws2b0n1_43, ws2b0n0_45, ws2b0n1_44, ws2b0n0_46, ws2b0n1_45, ws2b0n0_47, ws2b0n1_46, ws2b0n0_48, ws2b0n1_47, ws2b0n0_49, ws2b0n1_48, ws2b0n0_50, ws2b0n1_49, ws2b0n0_51, ws2b0n1_50, ws2b0n0_52, ws2b0n1_51, ws2b0n0_53, ws2b0n1_52, ws2b0n0_54, ws2b0n1_53, ws2b0n0_55, ws2b0n1_54, ws2b0n0_56, ws2b0n1_55, ws2b0n0_57, ws2b0n1_56, ws2b0n0_58, ws2b0n1_57, ws2b0n0_59, ws2b0n1_58, ws2b0n0_60, ws2b0n1_59, ws2b0n0_61, ws2b0n0_62, ws2b0n0_63, ws2b1n0_18, ws2b1n0_19, ws2b1n0_20, ws2b1n1_19, ws2b1n0_21, ws2b1n1_20, ws2b1n0_22, ws2b1n1_21, ws2b1n0_23, ws2b1n1_22, ws2b1n0_24, ws2b1n1_23, ws2b1n0_25, ws2b1n1_24, ws2b1n0_26, ws2b1n1_25, ws2b1n0_27, ws2b1n1_26, ws2b1n0_28, ws2b1n1_27, ws2b1n0_29, ws2b1n1_28, ws2b1n0_30, ws2b1n1_29, ws2b1n0_31, ws2b1n1_30, ws2b1n0_32, ws2b1n1_31, ws2b1n0_33, ws2b1n1_32, ws2b1n0_34, ws2b1n1_33, ws2b1n0_35, ws2b1n1_34, ws2b1n0_36, ws2b1n1_35, ws2b1n0_37, ws2b1n1_36, ws2b1n0_38, ws2b1n1_37, ws2b1n0_39, ws2b1n1_38, ws2b1n0_40, ws2b1n1_39, ws2b1n0_41, ws2b1n1_40, ws2b1n0_42, ws2b1n1_41, ws2b1n0_43, ws2b1n1_42, ws2b1n0_44, ws2b1n1_43, ws2b1n0_45, ws2b1n1_44, ws2b1n0_46, ws2b1n1_45, ws2b1n0_47, ws2b1n1_46, ws2b1n0_48, ws2b1n1_47, ws2b1n0_49, ws2b1n1_48, ws2b1n0_50, ws2b1n1_49, ws2b1n0_51, ws2b1n1_50, ws2b1n0_52, ws2b1n1_51, ws2b1n0_53, ws2b1n1_52, ws2b1n0_54, ws2b1n1_53, ws2b1n0_55, ws2b1n0_56, ws2b2n0_9, ws2b2n0_10, ws2b2n0_11, ws2b2n0_12, ws2b2n0_13, ws2b2n0_14, ws2b2n1_13, ws2b2n0_15, ws2b2n1_14, ws2b2n0_16, ws2b2n1_15, ws2b2n0_17, ws2b2n1_16, ws2b2n0_18, ws2b2n1_17, ws2b2n0_19, ws2b2n1_18, ws2b2n0_20, ws2b2n1_19, ws2b2n0_21, ws2b2n1_20, ws2b2n0_22, ws2b2n1_21, ws2b2n0_23, ws2b2n1_22, ws2b2n0_24, ws2b2n1_23, ws2b2n0_25, ws2b2n1_24, ws2b2n0_26, ws2b2n1_25, ws2b2n0_27, ws2b2n1_26, ws2b2n0_28, ws2b2n1_27, ws2b2n0_29, ws2b2n1_28, ws2b2n0_30, ws2b2n1_29, ws2b2n0_31, ws2b2n1_30, ws2b2n0_32, ws2b2n1_31, ws2b2n0_33, ws2b2n1_32, ws2b2n0_34, ws2b2n1_33, ws2b2n0_35, ws2b2n1_34, ws2b2n0_36, ws2b2n1_35, ws2b2n0_37, ws2b2n1_36, ws2b2n0_38, ws2b2n1_37, ws2b2n0_39, ws2b2n1_38, ws2b2n0_40, ws2b2n1_39, ws2b2n0_41, ws2b2n1_40, ws2b2n0_42, ws2b2n1_41, ws2b2n0_43, ws2b2n1_42, ws2b2n0_44, ws2b2n1_43, ws2b2n0_45, ws2b2n1_44, ws2b2n0_46, ws2b2n1_45, ws2b2n0_47, ws2b2n1_46, ws2b2n0_48, ws2b2n0_49, ws2b3n0_5, ws2b3n0_6, ws2b3n1_5, ws2b3n0_7, ws2b3n1_6, ws2b3n0_8, ws2b3n1_7, ws2b3n0_9, ws2b3n1_8, ws2b3n0_10, ws2b3n1_9, ws2b3n0_11, ws2b3n1_10, ws2b3n0_12, ws2b3n1_11, ws2b3n0_13, ws2b3n1_12, ws2b3n0_14, ws2b3n1_13, ws2b3n0_15, ws2b3n1_14, ws2b3n0_16, ws2b3n1_15, ws2b3n0_17, ws2b3n1_16, ws2b3n0_18, ws2b3n1_17, ws2b3n0_19, ws2b3n1_18, ws2b3n0_20, ws2b3n1_19, ws2b3n0_21, ws2b3n1_20, ws2b3n0_22, ws2b3n1_21, ws2b3n0_23, ws2b3n1_22, ws2b3n0_24, ws2b3n1_23, ws2b3n0_25, ws2b3n1_24, ws2b3n0_26, ws2b3n1_25, ws2b3n0_27, ws2b3n1_26, ws2b3n0_28, ws2b3n1_27, ws2b3n0_29, ws2b3n1_28, ws2b3n0_30, ws2b3n1_29, ws2b3n0_31, ws2b3n1_30, ws2b3n0_32, ws2b3n1_31, ws2b3n0_33, ws2b3n1_32, ws2b3n0_34, ws2b3n1_33, ws2b3n0_35, ws2b3n1_34, ws2b3n0_36, ws2b3n1_35, ws2b3n0_37, ws2b3n1_36, ws2b3n0_38, ws2b3n1_37, ws2b3n0_39, ws2b3n1_38, ws2b3n0_40, ws2b3n1_39, ws2b3n0_41, ws2b3n0_42, ws2b4n0_1, ws2b4n0_2, ws2b4n1_1, ws2b4n0_3, ws2b4n1_2, ws2b4n0_4, ws2b4n1_3, ws2b4n0_5, ws2b4n1_4, ws2b4n0_6, ws2b4n1_5, ws2b4n0_7, ws2b4n1_6, ws2b4n0_8, ws2b4n1_7, ws2b4n0_9, ws2b4n1_8, ws2b4n0_10, ws2b4n1_9, ws2b4n0_11, ws2b4n1_10, ws2b4n0_12, ws2b4n1_11, ws2b4n0_13, ws2b4n1_12, ws2b4n0_14, ws2b4n1_13, ws2b4n0_15, ws2b4n1_14, ws2b4n0_16, ws2b4n1_15, ws2b4n0_17, ws2b4n1_16, ws2b4n0_18, ws2b4n1_17, ws2b4n0_19, ws2b4n1_18, ws2b4n0_20, ws2b4n1_19, ws2b4n0_21, ws2b4n1_20, ws2b4n0_22, ws2b4n1_21, ws2b4n0_23, ws2b4n1_22, ws2b4n0_24, ws2b4n1_23, ws2b4n0_25, ws2b4n1_24, ws2b4n0_26, ws2b4n1_25, ws2b4n0_27, ws2b4n1_26, ws2b4n0_28, ws2b4n1_27, ws2b4n0_29, ws2b4n1_28, ws2b4n0_30, ws2b4n1_29, ws2b4n0_31, ws2b4n1_30, ws2b4n0_32, ws2b4n1_31, ws2b4n0_33, ws2b4n1_32, ws2b4n0_34, ws2b4n0_35, ws2b4n0_36;
wire ws3b0n0_18, ws3b0n0_19, ws3b0n0_20, ws3b0n0_21, ws3b0n0_22, ws3b0n0_23, ws3b0n0_24, ws3b0n1_23, ws3b0n0_25, ws3b0n1_24, ws3b0n0_26, ws3b0n1_25, ws3b0n0_27, ws3b0n1_26, ws3b0n0_28, ws3b0n1_27, ws3b0n0_29, ws3b0n1_28, ws3b0n0_30, ws3b0n1_29, ws3b0n0_31, ws3b0n1_30, ws3b0n0_32, ws3b0n1_31, ws3b0n0_33, ws3b0n1_32, ws3b0n0_34, ws3b0n1_33, ws3b0n0_35, ws3b0n1_34, ws3b0n0_36, ws3b0n1_35, ws3b0n0_37, ws3b0n1_36, ws3b0n0_38, ws3b0n1_37, ws3b0n0_39, ws3b0n1_38, ws3b0n0_40, ws3b0n1_39, ws3b0n0_41, ws3b0n1_40, ws3b0n0_42, ws3b0n1_41, ws3b0n0_43, ws3b0n1_42, ws3b0n0_44, ws3b0n1_43, ws3b0n0_45, ws3b0n1_44, ws3b0n0_46, ws3b0n1_45, ws3b0n0_47, ws3b0n1_46, ws3b0n0_48, ws3b0n1_47, ws3b0n0_49, ws3b0n1_48, ws3b0n0_50, ws3b0n1_49, ws3b0n0_51, ws3b0n1_50, ws3b0n0_52, ws3b0n1_51, ws3b0n0_53, ws3b0n1_52, ws3b0n0_54, ws3b0n1_53, ws3b0n0_55, ws3b0n1_54, ws3b0n0_56, ws3b0n1_55, ws3b0n0_57, ws3b0n1_56, ws3b0n0_58, ws3b0n1_57, ws3b0n0_59, ws3b0n1_58, ws3b0n0_60, ws3b0n0_61, ws3b0n0_62, ws3b0n0_63, ws3b1n0_9, ws3b1n0_10, ws3b1n0_11, ws3b1n0_12, ws3b1n0_13, ws3b1n1_12, ws3b1n0_14, ws3b1n1_13, ws3b1n0_15, ws3b1n1_14, ws3b1n0_16, ws3b1n1_15, ws3b1n0_17, ws3b1n1_16, ws3b1n0_18, ws3b1n1_17, ws3b1n0_19, ws3b1n1_18, ws3b1n0_20, ws3b1n1_19, ws3b1n0_21, ws3b1n1_20, ws3b1n0_22, ws3b1n1_21, ws3b1n0_23, ws3b1n1_22, ws3b1n0_24, ws3b1n1_23, ws3b1n0_25, ws3b1n1_24, ws3b1n0_26, ws3b1n1_25, ws3b1n0_27, ws3b1n1_26, ws3b1n0_28, ws3b1n1_27, ws3b1n0_29, ws3b1n1_28, ws3b1n0_30, ws3b1n1_29, ws3b1n0_31, ws3b1n1_30, ws3b1n0_32, ws3b1n1_31, ws3b1n0_33, ws3b1n1_32, ws3b1n0_34, ws3b1n1_33, ws3b1n0_35, ws3b1n1_34, ws3b1n0_36, ws3b1n1_35, ws3b1n0_37, ws3b1n1_36, ws3b1n0_38, ws3b1n1_37, ws3b1n0_39, ws3b1n1_38, ws3b1n0_40, ws3b1n1_39, ws3b1n0_41, ws3b1n1_40, ws3b1n0_42, ws3b1n1_41, ws3b1n0_43, ws3b1n1_42, ws3b1n0_44, ws3b1n1_43, ws3b1n0_45, ws3b1n1_44, ws3b1n0_46, ws3b1n1_45, ws3b1n0_47, ws3b1n1_46, ws3b1n0_48, ws3b1n1_47, ws3b1n0_49, ws3b1n1_48, ws3b1n0_50, ws3b1n0_51, ws3b1n0_52, ws3b1n0_53, ws3b2n0_1, ws3b2n0_2, ws3b2n0_3, ws3b2n0_4, ws3b2n0_5, ws3b2n1_4, ws3b2n0_6, ws3b2n1_5, ws3b2n0_7, ws3b2n1_6, ws3b2n0_8, ws3b2n1_7, ws3b2n0_9, ws3b2n1_8, ws3b2n0_10, ws3b2n1_9, ws3b2n0_11, ws3b2n1_10, ws3b2n0_12, ws3b2n1_11, ws3b2n0_13, ws3b2n1_12, ws3b2n0_14, ws3b2n1_13, ws3b2n0_15, ws3b2n1_14, ws3b2n0_16, ws3b2n1_15, ws3b2n0_17, ws3b2n1_16, ws3b2n0_18, ws3b2n1_17, ws3b2n0_19, ws3b2n1_18, ws3b2n0_20, ws3b2n1_19, ws3b2n0_21, ws3b2n1_20, ws3b2n0_22, ws3b2n1_21, ws3b2n0_23, ws3b2n1_22, ws3b2n0_24, ws3b2n1_23, ws3b2n0_25, ws3b2n1_24, ws3b2n0_26, ws3b2n1_25, ws3b2n0_27, ws3b2n1_26, ws3b2n0_28, ws3b2n1_27, ws3b2n0_29, ws3b2n1_28, ws3b2n0_30, ws3b2n1_29, ws3b2n0_31, ws3b2n1_30, ws3b2n0_32, ws3b2n1_31, ws3b2n0_33, ws3b2n1_32, ws3b2n0_34, ws3b2n1_33, ws3b2n0_35, ws3b2n1_34, ws3b2n0_36, ws3b2n1_35, ws3b2n0_37, ws3b2n1_36, ws3b2n0_38, ws3b2n1_37, ws3b2n0_39, ws3b2n1_38, ws3b2n0_40, ws3b2n0_41, ws3b2n0_42;
wire ws4b0n0_9, ws4b0n0_10, ws4b0n0_11, ws4b0n0_12, ws4b0n0_13, ws4b0n0_14, ws4b0n0_15, ws4b0n0_16, ws4b0n0_17, ws4b0n0_18, ws4b0n1_17, ws4b0n0_19, ws4b0n1_18, ws4b0n0_20, ws4b0n1_19, ws4b0n0_21, ws4b0n1_20, ws4b0n0_22, ws4b0n1_21, ws4b0n0_23, ws4b0n1_22, ws4b0n0_24, ws4b0n1_23, ws4b0n0_25, ws4b0n1_24, ws4b0n0_26, ws4b0n1_25, ws4b0n0_27, ws4b0n1_26, ws4b0n0_28, ws4b0n1_27, ws4b0n0_29, ws4b0n1_28, ws4b0n0_30, ws4b0n1_29, ws4b0n0_31, ws4b0n1_30, ws4b0n0_32, ws4b0n1_31, ws4b0n0_33, ws4b0n1_32, ws4b0n0_34, ws4b0n1_33, ws4b0n0_35, ws4b0n1_34, ws4b0n0_36, ws4b0n1_35, ws4b0n0_37, ws4b0n1_36, ws4b0n0_38, ws4b0n1_37, ws4b0n0_39, ws4b0n1_38, ws4b0n0_40, ws4b0n1_39, ws4b0n0_41, ws4b0n1_40, ws4b0n0_42, ws4b0n1_41, ws4b0n0_43, ws4b0n1_42, ws4b0n0_44, ws4b0n1_43, ws4b0n0_45, ws4b0n1_44, ws4b0n0_46, ws4b0n1_45, ws4b0n0_47, ws4b0n1_46, ws4b0n0_48, ws4b0n1_47, ws4b0n0_49, ws4b0n1_48, ws4b0n0_50, ws4b0n1_49, ws4b0n0_51, ws4b0n1_50, ws4b0n0_52, ws4b0n1_51, ws4b0n0_53, ws4b0n1_52, ws4b0n0_54, ws4b0n1_53, ws4b0n0_55, ws4b0n1_54, ws4b0n0_56, ws4b0n1_55, ws4b0n0_57, ws4b0n1_56, ws4b0n0_58, ws4b0n1_57, ws4b0n0_59, ws4b0n0_60, ws4b0n0_61, ws4b0n0_62, ws4b0n0_63, ws4b1n0_1, ws4b1n0_2, ws4b1n0_3, ws4b1n0_4, ws4b1n1_3, ws4b1n0_5, ws4b1n1_4, ws4b1n0_6, ws4b1n1_5, ws4b1n0_7, ws4b1n1_6, ws4b1n0_8, ws4b1n1_7, ws4b1n0_9, ws4b1n1_8, ws4b1n0_10, ws4b1n1_9, ws4b1n0_11, ws4b1n1_10, ws4b1n0_12, ws4b1n1_11, ws4b1n0_13, ws4b1n1_12, ws4b1n0_14, ws4b1n1_13, ws4b1n0_15, ws4b1n1_14, ws4b1n0_16, ws4b1n1_15, ws4b1n0_17, ws4b1n1_16, ws4b1n0_18, ws4b1n1_17, ws4b1n0_19, ws4b1n1_18, ws4b1n0_20, ws4b1n1_19, ws4b1n0_21, ws4b1n1_20, ws4b1n0_22, ws4b1n1_21, ws4b1n0_23, ws4b1n1_22, ws4b1n0_24, ws4b1n1_23, ws4b1n0_25, ws4b1n1_24, ws4b1n0_26, ws4b1n1_25, ws4b1n0_27, ws4b1n1_26, ws4b1n0_28, ws4b1n1_27, ws4b1n0_29, ws4b1n1_28, ws4b1n0_30, ws4b1n1_29, ws4b1n0_31, ws4b1n1_30, ws4b1n0_32, ws4b1n1_31, ws4b1n0_33, ws4b1n1_32, ws4b1n0_34, ws4b1n1_33, ws4b1n0_35, ws4b1n1_34, ws4b1n0_36, ws4b1n1_35, ws4b1n0_37, ws4b1n1_36, ws4b1n0_38, ws4b1n1_37, ws4b1n0_39, ws4b1n1_38, ws4b1n0_40, ws4b1n1_39, ws4b1n0_41, ws4b1n1_40, ws4b1n0_42, ws4b1n1_41, ws4b1n0_43, ws4b1n0_44, ws4b1n0_45, ws4b1n0_46, ws4b1n0_47, ws4b1n0_48;
wire ws5b0n0_1, ws5b0n0_2, ws5b0n0_3, ws5b0n0_4, ws5b0n0_5, ws5b0n0_6, ws5b0n0_7, ws5b0n0_8, ws5b0n0_9, ws5b0n1_8, ws5b0n0_10, ws5b0n1_9, ws5b0n0_11, ws5b0n1_10, ws5b0n0_12, ws5b0n1_11, ws5b0n0_13, ws5b0n1_12, ws5b0n0_14, ws5b0n1_13, ws5b0n0_15, ws5b0n1_14, ws5b0n0_16, ws5b0n1_15, ws5b0n0_17, ws5b0n1_16, ws5b0n0_18, ws5b0n1_17, ws5b0n0_19, ws5b0n1_18, ws5b0n0_20, ws5b0n1_19, ws5b0n0_21, ws5b0n1_20, ws5b0n0_22, ws5b0n1_21, ws5b0n0_23, ws5b0n1_22, ws5b0n0_24, ws5b0n1_23, ws5b0n0_25, ws5b0n1_24, ws5b0n0_26, ws5b0n1_25, ws5b0n0_27, ws5b0n1_26, ws5b0n0_28, ws5b0n1_27, ws5b0n0_29, ws5b0n1_28, ws5b0n0_30, ws5b0n1_29, ws5b0n0_31, ws5b0n1_30, ws5b0n0_32, ws5b0n1_31, ws5b0n0_33, ws5b0n1_32, ws5b0n0_34, ws5b0n1_33, ws5b0n0_35, ws5b0n1_34, ws5b0n0_36, ws5b0n1_35, ws5b0n0_37, ws5b0n1_36, ws5b0n0_38, ws5b0n1_37, ws5b0n0_39, ws5b0n1_38, ws5b0n0_40, ws5b0n1_39, ws5b0n0_41, ws5b0n1_40, ws5b0n0_42, ws5b0n1_41, ws5b0n0_43, ws5b0n1_42, ws5b0n0_44, ws5b0n1_43, ws5b0n0_45, ws5b0n1_44, ws5b0n0_46, ws5b0n1_45, ws5b0n0_47, ws5b0n1_46, ws5b0n0_48, ws5b0n1_47, ws5b0n0_49, ws5b0n1_48, ws5b0n0_50, ws5b0n1_49, ws5b0n0_51, ws5b0n1_50, ws5b0n0_52, ws5b0n1_51, ws5b0n0_53, ws5b0n1_52, ws5b0n0_54, ws5b0n1_53, ws5b0n0_55, ws5b0n1_54, ws5b0n0_56, ws5b0n1_55, ws5b0n0_57, ws5b0n1_56, ws5b0n0_58, ws5b0n0_59, ws5b0n0_60, ws5b0n0_61, ws5b0n0_62, ws5b0n0_63;
wire ws6b0n0_1, ws6b0n0_2, ws6b0n0_3, ws6b0n1_2, ws6b0n0_4, ws6b0n1_3, ws6b0n0_5, ws6b0n1_4, ws6b0n0_6, ws6b0n1_5, ws6b0n0_7, ws6b0n1_6, ws6b0n0_8, ws6b0n1_7, ws6b0n0_9, ws6b0n1_8, ws6b0n0_10, ws6b0n1_9, ws6b0n0_11, ws6b0n1_10, ws6b0n0_12, ws6b0n1_11, ws6b0n0_13, ws6b0n1_12, ws6b0n0_14, ws6b0n1_13, ws6b0n0_15, ws6b0n1_14, ws6b0n0_16, ws6b0n1_15, ws6b0n0_17, ws6b0n1_16, ws6b0n0_18, ws6b0n1_17, ws6b0n0_19, ws6b0n1_18, ws6b0n0_20, ws6b0n1_19, ws6b0n0_21, ws6b0n1_20, ws6b0n0_22, ws6b0n1_21, ws6b0n0_23, ws6b0n1_22, ws6b0n0_24, ws6b0n1_23, ws6b0n0_25, ws6b0n1_24, ws6b0n0_26, ws6b0n1_25, ws6b0n0_27, ws6b0n1_26, ws6b0n0_28, ws6b0n1_27, ws6b0n0_29, ws6b0n1_28, ws6b0n0_30, ws6b0n1_29, ws6b0n0_31, ws6b0n1_30, ws6b0n0_32, ws6b0n1_31, ws6b0n0_33, ws6b0n1_32, ws6b0n0_34, ws6b0n1_33, ws6b0n0_35, ws6b0n1_34, ws6b0n0_36, ws6b0n1_35, ws6b0n0_37, ws6b0n1_36, ws6b0n0_38, ws6b0n1_37, ws6b0n0_39, ws6b0n1_38, ws6b0n0_40, ws6b0n1_39, ws6b0n0_41, ws6b0n1_40, ws6b0n0_42, ws6b0n1_41, ws6b0n0_43, ws6b0n1_42, ws6b0n0_44, ws6b0n1_43, ws6b0n0_45, ws6b0n1_44, ws6b0n0_46, ws6b0n1_45, ws6b0n0_47, ws6b0n1_46, ws6b0n0_48, ws6b0n1_47, ws6b0n0_49, ws6b0n1_48, ws6b0n0_50, ws6b0n1_49, ws6b0n0_51, ws6b0n1_50, ws6b0n0_52, ws6b0n1_51, ws6b0n0_53, ws6b0n1_52, ws6b0n0_54, ws6b0n1_53, ws6b0n0_55, ws6b0n1_54, ws6b0n0_56, ws6b0n1_55, ws6b0n0_57, ws6b0n0_58, ws6b0n0_59, ws6b0n0_60, ws6b0n0_61, ws6b0n0_62, ws6b0n0_63;
wire ws7b0n0_1, ws7b0n1_0, ws7b0n0_2, ws7b0n1_1, ws7b0n0_3, ws7b0n1_2, ws7b0n0_4, ws7b0n1_3, ws7b0n0_5, ws7b0n1_4, ws7b0n0_6, ws7b0n1_5, ws7b0n0_7, ws7b0n1_6, ws7b0n0_8, ws7b0n1_7, ws7b0n0_9, ws7b0n1_8, ws7b0n0_10, ws7b0n1_9, ws7b0n0_11, ws7b0n1_10, ws7b0n0_12, ws7b0n1_11, ws7b0n0_13, ws7b0n1_12, ws7b0n0_14, ws7b0n1_13, ws7b0n0_15, ws7b0n1_14, ws7b0n0_16, ws7b0n1_15, ws7b0n0_17, ws7b0n1_16, ws7b0n0_18, ws7b0n1_17, ws7b0n0_19, ws7b0n1_18, ws7b0n0_20, ws7b0n1_19, ws7b0n0_21, ws7b0n1_20, ws7b0n0_22, ws7b0n1_21, ws7b0n0_23, ws7b0n1_22, ws7b0n0_24, ws7b0n1_23, ws7b0n0_25, ws7b0n1_24, ws7b0n0_26, ws7b0n1_25, ws7b0n0_27, ws7b0n1_26, ws7b0n0_28, ws7b0n1_27, ws7b0n0_29, ws7b0n1_28, ws7b0n0_30, ws7b0n1_29, ws7b0n0_31, ws7b0n1_30, ws7b0n0_32, ws7b0n1_31, ws7b0n0_33, ws7b0n1_32, ws7b0n0_34, ws7b0n1_33, ws7b0n0_35, ws7b0n1_34, ws7b0n0_36, ws7b0n1_35, ws7b0n0_37, ws7b0n1_36, ws7b0n0_38, ws7b0n1_37, ws7b0n0_39, ws7b0n1_38, ws7b0n0_40, ws7b0n1_39, ws7b0n0_41, ws7b0n1_40, ws7b0n0_42, ws7b0n1_41, ws7b0n0_43, ws7b0n1_42, ws7b0n0_44, ws7b0n1_43, ws7b0n0_45, ws7b0n1_44, ws7b0n0_46, ws7b0n1_45, ws7b0n0_47, ws7b0n1_46, ws7b0n0_48, ws7b0n1_47, ws7b0n0_49, ws7b0n1_48, ws7b0n0_50, ws7b0n1_49, ws7b0n0_51, ws7b0n1_50, ws7b0n0_52, ws7b0n1_51, ws7b0n0_53, ws7b0n1_52, ws7b0n0_54, ws7b0n1_53, ws7b0n0_55, ws7b0n1_54, ws7b0n0_56, ws7b0n0_57, ws7b0n0_58, ws7b0n0_59, ws7b0n0_60, ws7b0n0_61, ws7b0n0_62, ws7b0n0_63;

nand nand31_0(wand31_0, a[31], b[0]);
and and30_0(wand30_0, a[30], b[0]);
and and29_0(wand29_0, a[29], b[0]);
and and28_0(wand28_0, a[28], b[0]);
and and27_0(wand27_0, a[27], b[0]);
and and26_0(wand26_0, a[26], b[0]);
and and25_0(wand25_0, a[25], b[0]);
and and24_0(wand24_0, a[24], b[0]);
and and23_0(wand23_0, a[23], b[0]);
and and22_0(wand22_0, a[22], b[0]);
and and21_0(wand21_0, a[21], b[0]);
and and20_0(wand20_0, a[20], b[0]);
and and19_0(wand19_0, a[19], b[0]);
and and18_0(wand18_0, a[18], b[0]);
and and17_0(wand17_0, a[17], b[0]);
and and16_0(wand16_0, a[16], b[0]);
and and15_0(wand15_0, a[15], b[0]);
and and14_0(wand14_0, a[14], b[0]);
and and13_0(wand13_0, a[13], b[0]);
and and12_0(wand12_0, a[12], b[0]);
and and11_0(wand11_0, a[11], b[0]);
and and10_0(wand10_0, a[10], b[0]);
and and9_0(wand9_0, a[9], b[0]);
and and8_0(wand8_0, a[8], b[0]);
and and7_0(wand7_0, a[7], b[0]);
and and6_0(wand6_0, a[6], b[0]);
and and5_0(wand5_0, a[5], b[0]);
and and4_0(wand4_0, a[4], b[0]);
and and3_0(wand3_0, a[3], b[0]);
and and2_0(wand2_0, a[2], b[0]);
and and1_0(wand1_0, a[1], b[0]);
and and0_0(wand0_0, a[0], b[0]);
nand nand31_1(wand31_1, a[31], b[1]);
and and30_1(wand30_1, a[30], b[1]);
and and29_1(wand29_1, a[29], b[1]);
and and28_1(wand28_1, a[28], b[1]);
and and27_1(wand27_1, a[27], b[1]);
and and26_1(wand26_1, a[26], b[1]);
and and25_1(wand25_1, a[25], b[1]);
and and24_1(wand24_1, a[24], b[1]);
and and23_1(wand23_1, a[23], b[1]);
and and22_1(wand22_1, a[22], b[1]);
and and21_1(wand21_1, a[21], b[1]);
and and20_1(wand20_1, a[20], b[1]);
and and19_1(wand19_1, a[19], b[1]);
and and18_1(wand18_1, a[18], b[1]);
and and17_1(wand17_1, a[17], b[1]);
and and16_1(wand16_1, a[16], b[1]);
and and15_1(wand15_1, a[15], b[1]);
and and14_1(wand14_1, a[14], b[1]);
and and13_1(wand13_1, a[13], b[1]);
and and12_1(wand12_1, a[12], b[1]);
and and11_1(wand11_1, a[11], b[1]);
and and10_1(wand10_1, a[10], b[1]);
and and9_1(wand9_1, a[9], b[1]);
and and8_1(wand8_1, a[8], b[1]);
and and7_1(wand7_1, a[7], b[1]);
and and6_1(wand6_1, a[6], b[1]);
and and5_1(wand5_1, a[5], b[1]);
and and4_1(wand4_1, a[4], b[1]);
and and3_1(wand3_1, a[3], b[1]);
and and2_1(wand2_1, a[2], b[1]);
and and1_1(wand1_1, a[1], b[1]);
and and0_1(wand0_1, a[0], b[1]);
nand nand31_2(wand31_2, a[31], b[2]);
and and30_2(wand30_2, a[30], b[2]);
and and29_2(wand29_2, a[29], b[2]);
and and28_2(wand28_2, a[28], b[2]);
and and27_2(wand27_2, a[27], b[2]);
and and26_2(wand26_2, a[26], b[2]);
and and25_2(wand25_2, a[25], b[2]);
and and24_2(wand24_2, a[24], b[2]);
and and23_2(wand23_2, a[23], b[2]);
and and22_2(wand22_2, a[22], b[2]);
and and21_2(wand21_2, a[21], b[2]);
and and20_2(wand20_2, a[20], b[2]);
and and19_2(wand19_2, a[19], b[2]);
and and18_2(wand18_2, a[18], b[2]);
and and17_2(wand17_2, a[17], b[2]);
and and16_2(wand16_2, a[16], b[2]);
and and15_2(wand15_2, a[15], b[2]);
and and14_2(wand14_2, a[14], b[2]);
and and13_2(wand13_2, a[13], b[2]);
and and12_2(wand12_2, a[12], b[2]);
and and11_2(wand11_2, a[11], b[2]);
and and10_2(wand10_2, a[10], b[2]);
and and9_2(wand9_2, a[9], b[2]);
and and8_2(wand8_2, a[8], b[2]);
and and7_2(wand7_2, a[7], b[2]);
and and6_2(wand6_2, a[6], b[2]);
and and5_2(wand5_2, a[5], b[2]);
and and4_2(wand4_2, a[4], b[2]);
and and3_2(wand3_2, a[3], b[2]);
and and2_2(wand2_2, a[2], b[2]);
and and1_2(wand1_2, a[1], b[2]);
and and0_2(wand0_2, a[0], b[2]);
nand nand31_3(wand31_3, a[31], b[3]);
and and30_3(wand30_3, a[30], b[3]);
and and29_3(wand29_3, a[29], b[3]);
and and28_3(wand28_3, a[28], b[3]);
and and27_3(wand27_3, a[27], b[3]);
and and26_3(wand26_3, a[26], b[3]);
and and25_3(wand25_3, a[25], b[3]);
and and24_3(wand24_3, a[24], b[3]);
and and23_3(wand23_3, a[23], b[3]);
and and22_3(wand22_3, a[22], b[3]);
and and21_3(wand21_3, a[21], b[3]);
and and20_3(wand20_3, a[20], b[3]);
and and19_3(wand19_3, a[19], b[3]);
and and18_3(wand18_3, a[18], b[3]);
and and17_3(wand17_3, a[17], b[3]);
and and16_3(wand16_3, a[16], b[3]);
and and15_3(wand15_3, a[15], b[3]);
and and14_3(wand14_3, a[14], b[3]);
and and13_3(wand13_3, a[13], b[3]);
and and12_3(wand12_3, a[12], b[3]);
and and11_3(wand11_3, a[11], b[3]);
and and10_3(wand10_3, a[10], b[3]);
and and9_3(wand9_3, a[9], b[3]);
and and8_3(wand8_3, a[8], b[3]);
and and7_3(wand7_3, a[7], b[3]);
and and6_3(wand6_3, a[6], b[3]);
and and5_3(wand5_3, a[5], b[3]);
and and4_3(wand4_3, a[4], b[3]);
and and3_3(wand3_3, a[3], b[3]);
and and2_3(wand2_3, a[2], b[3]);
and and1_3(wand1_3, a[1], b[3]);
and and0_3(wand0_3, a[0], b[3]);
nand nand31_4(wand31_4, a[31], b[4]);
and and30_4(wand30_4, a[30], b[4]);
and and29_4(wand29_4, a[29], b[4]);
and and28_4(wand28_4, a[28], b[4]);
and and27_4(wand27_4, a[27], b[4]);
and and26_4(wand26_4, a[26], b[4]);
and and25_4(wand25_4, a[25], b[4]);
and and24_4(wand24_4, a[24], b[4]);
and and23_4(wand23_4, a[23], b[4]);
and and22_4(wand22_4, a[22], b[4]);
and and21_4(wand21_4, a[21], b[4]);
and and20_4(wand20_4, a[20], b[4]);
and and19_4(wand19_4, a[19], b[4]);
and and18_4(wand18_4, a[18], b[4]);
and and17_4(wand17_4, a[17], b[4]);
and and16_4(wand16_4, a[16], b[4]);
and and15_4(wand15_4, a[15], b[4]);
and and14_4(wand14_4, a[14], b[4]);
and and13_4(wand13_4, a[13], b[4]);
and and12_4(wand12_4, a[12], b[4]);
and and11_4(wand11_4, a[11], b[4]);
and and10_4(wand10_4, a[10], b[4]);
and and9_4(wand9_4, a[9], b[4]);
and and8_4(wand8_4, a[8], b[4]);
and and7_4(wand7_4, a[7], b[4]);
and and6_4(wand6_4, a[6], b[4]);
and and5_4(wand5_4, a[5], b[4]);
and and4_4(wand4_4, a[4], b[4]);
and and3_4(wand3_4, a[3], b[4]);
and and2_4(wand2_4, a[2], b[4]);
and and1_4(wand1_4, a[1], b[4]);
and and0_4(wand0_4, a[0], b[4]);
nand nand31_5(wand31_5, a[31], b[5]);
and and30_5(wand30_5, a[30], b[5]);
and and29_5(wand29_5, a[29], b[5]);
and and28_5(wand28_5, a[28], b[5]);
and and27_5(wand27_5, a[27], b[5]);
and and26_5(wand26_5, a[26], b[5]);
and and25_5(wand25_5, a[25], b[5]);
and and24_5(wand24_5, a[24], b[5]);
and and23_5(wand23_5, a[23], b[5]);
and and22_5(wand22_5, a[22], b[5]);
and and21_5(wand21_5, a[21], b[5]);
and and20_5(wand20_5, a[20], b[5]);
and and19_5(wand19_5, a[19], b[5]);
and and18_5(wand18_5, a[18], b[5]);
and and17_5(wand17_5, a[17], b[5]);
and and16_5(wand16_5, a[16], b[5]);
and and15_5(wand15_5, a[15], b[5]);
and and14_5(wand14_5, a[14], b[5]);
and and13_5(wand13_5, a[13], b[5]);
and and12_5(wand12_5, a[12], b[5]);
and and11_5(wand11_5, a[11], b[5]);
and and10_5(wand10_5, a[10], b[5]);
and and9_5(wand9_5, a[9], b[5]);
and and8_5(wand8_5, a[8], b[5]);
and and7_5(wand7_5, a[7], b[5]);
and and6_5(wand6_5, a[6], b[5]);
and and5_5(wand5_5, a[5], b[5]);
and and4_5(wand4_5, a[4], b[5]);
and and3_5(wand3_5, a[3], b[5]);
and and2_5(wand2_5, a[2], b[5]);
and and1_5(wand1_5, a[1], b[5]);
and and0_5(wand0_5, a[0], b[5]);
nand nand31_6(wand31_6, a[31], b[6]);
and and30_6(wand30_6, a[30], b[6]);
and and29_6(wand29_6, a[29], b[6]);
and and28_6(wand28_6, a[28], b[6]);
and and27_6(wand27_6, a[27], b[6]);
and and26_6(wand26_6, a[26], b[6]);
and and25_6(wand25_6, a[25], b[6]);
and and24_6(wand24_6, a[24], b[6]);
and and23_6(wand23_6, a[23], b[6]);
and and22_6(wand22_6, a[22], b[6]);
and and21_6(wand21_6, a[21], b[6]);
and and20_6(wand20_6, a[20], b[6]);
and and19_6(wand19_6, a[19], b[6]);
and and18_6(wand18_6, a[18], b[6]);
and and17_6(wand17_6, a[17], b[6]);
and and16_6(wand16_6, a[16], b[6]);
and and15_6(wand15_6, a[15], b[6]);
and and14_6(wand14_6, a[14], b[6]);
and and13_6(wand13_6, a[13], b[6]);
and and12_6(wand12_6, a[12], b[6]);
and and11_6(wand11_6, a[11], b[6]);
and and10_6(wand10_6, a[10], b[6]);
and and9_6(wand9_6, a[9], b[6]);
and and8_6(wand8_6, a[8], b[6]);
and and7_6(wand7_6, a[7], b[6]);
and and6_6(wand6_6, a[6], b[6]);
and and5_6(wand5_6, a[5], b[6]);
and and4_6(wand4_6, a[4], b[6]);
and and3_6(wand3_6, a[3], b[6]);
and and2_6(wand2_6, a[2], b[6]);
and and1_6(wand1_6, a[1], b[6]);
and and0_6(wand0_6, a[0], b[6]);
nand nand31_7(wand31_7, a[31], b[7]);
and and30_7(wand30_7, a[30], b[7]);
and and29_7(wand29_7, a[29], b[7]);
and and28_7(wand28_7, a[28], b[7]);
and and27_7(wand27_7, a[27], b[7]);
and and26_7(wand26_7, a[26], b[7]);
and and25_7(wand25_7, a[25], b[7]);
and and24_7(wand24_7, a[24], b[7]);
and and23_7(wand23_7, a[23], b[7]);
and and22_7(wand22_7, a[22], b[7]);
and and21_7(wand21_7, a[21], b[7]);
and and20_7(wand20_7, a[20], b[7]);
and and19_7(wand19_7, a[19], b[7]);
and and18_7(wand18_7, a[18], b[7]);
and and17_7(wand17_7, a[17], b[7]);
and and16_7(wand16_7, a[16], b[7]);
and and15_7(wand15_7, a[15], b[7]);
and and14_7(wand14_7, a[14], b[7]);
and and13_7(wand13_7, a[13], b[7]);
and and12_7(wand12_7, a[12], b[7]);
and and11_7(wand11_7, a[11], b[7]);
and and10_7(wand10_7, a[10], b[7]);
and and9_7(wand9_7, a[9], b[7]);
and and8_7(wand8_7, a[8], b[7]);
and and7_7(wand7_7, a[7], b[7]);
and and6_7(wand6_7, a[6], b[7]);
and and5_7(wand5_7, a[5], b[7]);
and and4_7(wand4_7, a[4], b[7]);
and and3_7(wand3_7, a[3], b[7]);
and and2_7(wand2_7, a[2], b[7]);
and and1_7(wand1_7, a[1], b[7]);
and and0_7(wand0_7, a[0], b[7]);
nand nand31_8(wand31_8, a[31], b[8]);
and and30_8(wand30_8, a[30], b[8]);
and and29_8(wand29_8, a[29], b[8]);
and and28_8(wand28_8, a[28], b[8]);
and and27_8(wand27_8, a[27], b[8]);
and and26_8(wand26_8, a[26], b[8]);
and and25_8(wand25_8, a[25], b[8]);
and and24_8(wand24_8, a[24], b[8]);
and and23_8(wand23_8, a[23], b[8]);
and and22_8(wand22_8, a[22], b[8]);
and and21_8(wand21_8, a[21], b[8]);
and and20_8(wand20_8, a[20], b[8]);
and and19_8(wand19_8, a[19], b[8]);
and and18_8(wand18_8, a[18], b[8]);
and and17_8(wand17_8, a[17], b[8]);
and and16_8(wand16_8, a[16], b[8]);
and and15_8(wand15_8, a[15], b[8]);
and and14_8(wand14_8, a[14], b[8]);
and and13_8(wand13_8, a[13], b[8]);
and and12_8(wand12_8, a[12], b[8]);
and and11_8(wand11_8, a[11], b[8]);
and and10_8(wand10_8, a[10], b[8]);
and and9_8(wand9_8, a[9], b[8]);
and and8_8(wand8_8, a[8], b[8]);
and and7_8(wand7_8, a[7], b[8]);
and and6_8(wand6_8, a[6], b[8]);
and and5_8(wand5_8, a[5], b[8]);
and and4_8(wand4_8, a[4], b[8]);
and and3_8(wand3_8, a[3], b[8]);
and and2_8(wand2_8, a[2], b[8]);
and and1_8(wand1_8, a[1], b[8]);
and and0_8(wand0_8, a[0], b[8]);
nand nand31_9(wand31_9, a[31], b[9]);
and and30_9(wand30_9, a[30], b[9]);
and and29_9(wand29_9, a[29], b[9]);
and and28_9(wand28_9, a[28], b[9]);
and and27_9(wand27_9, a[27], b[9]);
and and26_9(wand26_9, a[26], b[9]);
and and25_9(wand25_9, a[25], b[9]);
and and24_9(wand24_9, a[24], b[9]);
and and23_9(wand23_9, a[23], b[9]);
and and22_9(wand22_9, a[22], b[9]);
and and21_9(wand21_9, a[21], b[9]);
and and20_9(wand20_9, a[20], b[9]);
and and19_9(wand19_9, a[19], b[9]);
and and18_9(wand18_9, a[18], b[9]);
and and17_9(wand17_9, a[17], b[9]);
and and16_9(wand16_9, a[16], b[9]);
and and15_9(wand15_9, a[15], b[9]);
and and14_9(wand14_9, a[14], b[9]);
and and13_9(wand13_9, a[13], b[9]);
and and12_9(wand12_9, a[12], b[9]);
and and11_9(wand11_9, a[11], b[9]);
and and10_9(wand10_9, a[10], b[9]);
and and9_9(wand9_9, a[9], b[9]);
and and8_9(wand8_9, a[8], b[9]);
and and7_9(wand7_9, a[7], b[9]);
and and6_9(wand6_9, a[6], b[9]);
and and5_9(wand5_9, a[5], b[9]);
and and4_9(wand4_9, a[4], b[9]);
and and3_9(wand3_9, a[3], b[9]);
and and2_9(wand2_9, a[2], b[9]);
and and1_9(wand1_9, a[1], b[9]);
and and0_9(wand0_9, a[0], b[9]);
nand nand31_10(wand31_10, a[31], b[10]);
and and30_10(wand30_10, a[30], b[10]);
and and29_10(wand29_10, a[29], b[10]);
and and28_10(wand28_10, a[28], b[10]);
and and27_10(wand27_10, a[27], b[10]);
and and26_10(wand26_10, a[26], b[10]);
and and25_10(wand25_10, a[25], b[10]);
and and24_10(wand24_10, a[24], b[10]);
and and23_10(wand23_10, a[23], b[10]);
and and22_10(wand22_10, a[22], b[10]);
and and21_10(wand21_10, a[21], b[10]);
and and20_10(wand20_10, a[20], b[10]);
and and19_10(wand19_10, a[19], b[10]);
and and18_10(wand18_10, a[18], b[10]);
and and17_10(wand17_10, a[17], b[10]);
and and16_10(wand16_10, a[16], b[10]);
and and15_10(wand15_10, a[15], b[10]);
and and14_10(wand14_10, a[14], b[10]);
and and13_10(wand13_10, a[13], b[10]);
and and12_10(wand12_10, a[12], b[10]);
and and11_10(wand11_10, a[11], b[10]);
and and10_10(wand10_10, a[10], b[10]);
and and9_10(wand9_10, a[9], b[10]);
and and8_10(wand8_10, a[8], b[10]);
and and7_10(wand7_10, a[7], b[10]);
and and6_10(wand6_10, a[6], b[10]);
and and5_10(wand5_10, a[5], b[10]);
and and4_10(wand4_10, a[4], b[10]);
and and3_10(wand3_10, a[3], b[10]);
and and2_10(wand2_10, a[2], b[10]);
and and1_10(wand1_10, a[1], b[10]);
and and0_10(wand0_10, a[0], b[10]);
nand nand31_11(wand31_11, a[31], b[11]);
and and30_11(wand30_11, a[30], b[11]);
and and29_11(wand29_11, a[29], b[11]);
and and28_11(wand28_11, a[28], b[11]);
and and27_11(wand27_11, a[27], b[11]);
and and26_11(wand26_11, a[26], b[11]);
and and25_11(wand25_11, a[25], b[11]);
and and24_11(wand24_11, a[24], b[11]);
and and23_11(wand23_11, a[23], b[11]);
and and22_11(wand22_11, a[22], b[11]);
and and21_11(wand21_11, a[21], b[11]);
and and20_11(wand20_11, a[20], b[11]);
and and19_11(wand19_11, a[19], b[11]);
and and18_11(wand18_11, a[18], b[11]);
and and17_11(wand17_11, a[17], b[11]);
and and16_11(wand16_11, a[16], b[11]);
and and15_11(wand15_11, a[15], b[11]);
and and14_11(wand14_11, a[14], b[11]);
and and13_11(wand13_11, a[13], b[11]);
and and12_11(wand12_11, a[12], b[11]);
and and11_11(wand11_11, a[11], b[11]);
and and10_11(wand10_11, a[10], b[11]);
and and9_11(wand9_11, a[9], b[11]);
and and8_11(wand8_11, a[8], b[11]);
and and7_11(wand7_11, a[7], b[11]);
and and6_11(wand6_11, a[6], b[11]);
and and5_11(wand5_11, a[5], b[11]);
and and4_11(wand4_11, a[4], b[11]);
and and3_11(wand3_11, a[3], b[11]);
and and2_11(wand2_11, a[2], b[11]);
and and1_11(wand1_11, a[1], b[11]);
and and0_11(wand0_11, a[0], b[11]);
nand nand31_12(wand31_12, a[31], b[12]);
and and30_12(wand30_12, a[30], b[12]);
and and29_12(wand29_12, a[29], b[12]);
and and28_12(wand28_12, a[28], b[12]);
and and27_12(wand27_12, a[27], b[12]);
and and26_12(wand26_12, a[26], b[12]);
and and25_12(wand25_12, a[25], b[12]);
and and24_12(wand24_12, a[24], b[12]);
and and23_12(wand23_12, a[23], b[12]);
and and22_12(wand22_12, a[22], b[12]);
and and21_12(wand21_12, a[21], b[12]);
and and20_12(wand20_12, a[20], b[12]);
and and19_12(wand19_12, a[19], b[12]);
and and18_12(wand18_12, a[18], b[12]);
and and17_12(wand17_12, a[17], b[12]);
and and16_12(wand16_12, a[16], b[12]);
and and15_12(wand15_12, a[15], b[12]);
and and14_12(wand14_12, a[14], b[12]);
and and13_12(wand13_12, a[13], b[12]);
and and12_12(wand12_12, a[12], b[12]);
and and11_12(wand11_12, a[11], b[12]);
and and10_12(wand10_12, a[10], b[12]);
and and9_12(wand9_12, a[9], b[12]);
and and8_12(wand8_12, a[8], b[12]);
and and7_12(wand7_12, a[7], b[12]);
and and6_12(wand6_12, a[6], b[12]);
and and5_12(wand5_12, a[5], b[12]);
and and4_12(wand4_12, a[4], b[12]);
and and3_12(wand3_12, a[3], b[12]);
and and2_12(wand2_12, a[2], b[12]);
and and1_12(wand1_12, a[1], b[12]);
and and0_12(wand0_12, a[0], b[12]);
nand nand31_13(wand31_13, a[31], b[13]);
and and30_13(wand30_13, a[30], b[13]);
and and29_13(wand29_13, a[29], b[13]);
and and28_13(wand28_13, a[28], b[13]);
and and27_13(wand27_13, a[27], b[13]);
and and26_13(wand26_13, a[26], b[13]);
and and25_13(wand25_13, a[25], b[13]);
and and24_13(wand24_13, a[24], b[13]);
and and23_13(wand23_13, a[23], b[13]);
and and22_13(wand22_13, a[22], b[13]);
and and21_13(wand21_13, a[21], b[13]);
and and20_13(wand20_13, a[20], b[13]);
and and19_13(wand19_13, a[19], b[13]);
and and18_13(wand18_13, a[18], b[13]);
and and17_13(wand17_13, a[17], b[13]);
and and16_13(wand16_13, a[16], b[13]);
and and15_13(wand15_13, a[15], b[13]);
and and14_13(wand14_13, a[14], b[13]);
and and13_13(wand13_13, a[13], b[13]);
and and12_13(wand12_13, a[12], b[13]);
and and11_13(wand11_13, a[11], b[13]);
and and10_13(wand10_13, a[10], b[13]);
and and9_13(wand9_13, a[9], b[13]);
and and8_13(wand8_13, a[8], b[13]);
and and7_13(wand7_13, a[7], b[13]);
and and6_13(wand6_13, a[6], b[13]);
and and5_13(wand5_13, a[5], b[13]);
and and4_13(wand4_13, a[4], b[13]);
and and3_13(wand3_13, a[3], b[13]);
and and2_13(wand2_13, a[2], b[13]);
and and1_13(wand1_13, a[1], b[13]);
and and0_13(wand0_13, a[0], b[13]);
nand nand31_14(wand31_14, a[31], b[14]);
and and30_14(wand30_14, a[30], b[14]);
and and29_14(wand29_14, a[29], b[14]);
and and28_14(wand28_14, a[28], b[14]);
and and27_14(wand27_14, a[27], b[14]);
and and26_14(wand26_14, a[26], b[14]);
and and25_14(wand25_14, a[25], b[14]);
and and24_14(wand24_14, a[24], b[14]);
and and23_14(wand23_14, a[23], b[14]);
and and22_14(wand22_14, a[22], b[14]);
and and21_14(wand21_14, a[21], b[14]);
and and20_14(wand20_14, a[20], b[14]);
and and19_14(wand19_14, a[19], b[14]);
and and18_14(wand18_14, a[18], b[14]);
and and17_14(wand17_14, a[17], b[14]);
and and16_14(wand16_14, a[16], b[14]);
and and15_14(wand15_14, a[15], b[14]);
and and14_14(wand14_14, a[14], b[14]);
and and13_14(wand13_14, a[13], b[14]);
and and12_14(wand12_14, a[12], b[14]);
and and11_14(wand11_14, a[11], b[14]);
and and10_14(wand10_14, a[10], b[14]);
and and9_14(wand9_14, a[9], b[14]);
and and8_14(wand8_14, a[8], b[14]);
and and7_14(wand7_14, a[7], b[14]);
and and6_14(wand6_14, a[6], b[14]);
and and5_14(wand5_14, a[5], b[14]);
and and4_14(wand4_14, a[4], b[14]);
and and3_14(wand3_14, a[3], b[14]);
and and2_14(wand2_14, a[2], b[14]);
and and1_14(wand1_14, a[1], b[14]);
and and0_14(wand0_14, a[0], b[14]);
nand nand31_15(wand31_15, a[31], b[15]);
and and30_15(wand30_15, a[30], b[15]);
and and29_15(wand29_15, a[29], b[15]);
and and28_15(wand28_15, a[28], b[15]);
and and27_15(wand27_15, a[27], b[15]);
and and26_15(wand26_15, a[26], b[15]);
and and25_15(wand25_15, a[25], b[15]);
and and24_15(wand24_15, a[24], b[15]);
and and23_15(wand23_15, a[23], b[15]);
and and22_15(wand22_15, a[22], b[15]);
and and21_15(wand21_15, a[21], b[15]);
and and20_15(wand20_15, a[20], b[15]);
and and19_15(wand19_15, a[19], b[15]);
and and18_15(wand18_15, a[18], b[15]);
and and17_15(wand17_15, a[17], b[15]);
and and16_15(wand16_15, a[16], b[15]);
and and15_15(wand15_15, a[15], b[15]);
and and14_15(wand14_15, a[14], b[15]);
and and13_15(wand13_15, a[13], b[15]);
and and12_15(wand12_15, a[12], b[15]);
and and11_15(wand11_15, a[11], b[15]);
and and10_15(wand10_15, a[10], b[15]);
and and9_15(wand9_15, a[9], b[15]);
and and8_15(wand8_15, a[8], b[15]);
and and7_15(wand7_15, a[7], b[15]);
and and6_15(wand6_15, a[6], b[15]);
and and5_15(wand5_15, a[5], b[15]);
and and4_15(wand4_15, a[4], b[15]);
and and3_15(wand3_15, a[3], b[15]);
and and2_15(wand2_15, a[2], b[15]);
and and1_15(wand1_15, a[1], b[15]);
and and0_15(wand0_15, a[0], b[15]);
nand nand31_16(wand31_16, a[31], b[16]);
and and30_16(wand30_16, a[30], b[16]);
and and29_16(wand29_16, a[29], b[16]);
and and28_16(wand28_16, a[28], b[16]);
and and27_16(wand27_16, a[27], b[16]);
and and26_16(wand26_16, a[26], b[16]);
and and25_16(wand25_16, a[25], b[16]);
and and24_16(wand24_16, a[24], b[16]);
and and23_16(wand23_16, a[23], b[16]);
and and22_16(wand22_16, a[22], b[16]);
and and21_16(wand21_16, a[21], b[16]);
and and20_16(wand20_16, a[20], b[16]);
and and19_16(wand19_16, a[19], b[16]);
and and18_16(wand18_16, a[18], b[16]);
and and17_16(wand17_16, a[17], b[16]);
and and16_16(wand16_16, a[16], b[16]);
and and15_16(wand15_16, a[15], b[16]);
and and14_16(wand14_16, a[14], b[16]);
and and13_16(wand13_16, a[13], b[16]);
and and12_16(wand12_16, a[12], b[16]);
and and11_16(wand11_16, a[11], b[16]);
and and10_16(wand10_16, a[10], b[16]);
and and9_16(wand9_16, a[9], b[16]);
and and8_16(wand8_16, a[8], b[16]);
and and7_16(wand7_16, a[7], b[16]);
and and6_16(wand6_16, a[6], b[16]);
and and5_16(wand5_16, a[5], b[16]);
and and4_16(wand4_16, a[4], b[16]);
and and3_16(wand3_16, a[3], b[16]);
and and2_16(wand2_16, a[2], b[16]);
and and1_16(wand1_16, a[1], b[16]);
and and0_16(wand0_16, a[0], b[16]);
nand nand31_17(wand31_17, a[31], b[17]);
and and30_17(wand30_17, a[30], b[17]);
and and29_17(wand29_17, a[29], b[17]);
and and28_17(wand28_17, a[28], b[17]);
and and27_17(wand27_17, a[27], b[17]);
and and26_17(wand26_17, a[26], b[17]);
and and25_17(wand25_17, a[25], b[17]);
and and24_17(wand24_17, a[24], b[17]);
and and23_17(wand23_17, a[23], b[17]);
and and22_17(wand22_17, a[22], b[17]);
and and21_17(wand21_17, a[21], b[17]);
and and20_17(wand20_17, a[20], b[17]);
and and19_17(wand19_17, a[19], b[17]);
and and18_17(wand18_17, a[18], b[17]);
and and17_17(wand17_17, a[17], b[17]);
and and16_17(wand16_17, a[16], b[17]);
and and15_17(wand15_17, a[15], b[17]);
and and14_17(wand14_17, a[14], b[17]);
and and13_17(wand13_17, a[13], b[17]);
and and12_17(wand12_17, a[12], b[17]);
and and11_17(wand11_17, a[11], b[17]);
and and10_17(wand10_17, a[10], b[17]);
and and9_17(wand9_17, a[9], b[17]);
and and8_17(wand8_17, a[8], b[17]);
and and7_17(wand7_17, a[7], b[17]);
and and6_17(wand6_17, a[6], b[17]);
and and5_17(wand5_17, a[5], b[17]);
and and4_17(wand4_17, a[4], b[17]);
and and3_17(wand3_17, a[3], b[17]);
and and2_17(wand2_17, a[2], b[17]);
and and1_17(wand1_17, a[1], b[17]);
and and0_17(wand0_17, a[0], b[17]);
nand nand31_18(wand31_18, a[31], b[18]);
and and30_18(wand30_18, a[30], b[18]);
and and29_18(wand29_18, a[29], b[18]);
and and28_18(wand28_18, a[28], b[18]);
and and27_18(wand27_18, a[27], b[18]);
and and26_18(wand26_18, a[26], b[18]);
and and25_18(wand25_18, a[25], b[18]);
and and24_18(wand24_18, a[24], b[18]);
and and23_18(wand23_18, a[23], b[18]);
and and22_18(wand22_18, a[22], b[18]);
and and21_18(wand21_18, a[21], b[18]);
and and20_18(wand20_18, a[20], b[18]);
and and19_18(wand19_18, a[19], b[18]);
and and18_18(wand18_18, a[18], b[18]);
and and17_18(wand17_18, a[17], b[18]);
and and16_18(wand16_18, a[16], b[18]);
and and15_18(wand15_18, a[15], b[18]);
and and14_18(wand14_18, a[14], b[18]);
and and13_18(wand13_18, a[13], b[18]);
and and12_18(wand12_18, a[12], b[18]);
and and11_18(wand11_18, a[11], b[18]);
and and10_18(wand10_18, a[10], b[18]);
and and9_18(wand9_18, a[9], b[18]);
and and8_18(wand8_18, a[8], b[18]);
and and7_18(wand7_18, a[7], b[18]);
and and6_18(wand6_18, a[6], b[18]);
and and5_18(wand5_18, a[5], b[18]);
and and4_18(wand4_18, a[4], b[18]);
and and3_18(wand3_18, a[3], b[18]);
and and2_18(wand2_18, a[2], b[18]);
and and1_18(wand1_18, a[1], b[18]);
and and0_18(wand0_18, a[0], b[18]);
nand nand31_19(wand31_19, a[31], b[19]);
and and30_19(wand30_19, a[30], b[19]);
and and29_19(wand29_19, a[29], b[19]);
and and28_19(wand28_19, a[28], b[19]);
and and27_19(wand27_19, a[27], b[19]);
and and26_19(wand26_19, a[26], b[19]);
and and25_19(wand25_19, a[25], b[19]);
and and24_19(wand24_19, a[24], b[19]);
and and23_19(wand23_19, a[23], b[19]);
and and22_19(wand22_19, a[22], b[19]);
and and21_19(wand21_19, a[21], b[19]);
and and20_19(wand20_19, a[20], b[19]);
and and19_19(wand19_19, a[19], b[19]);
and and18_19(wand18_19, a[18], b[19]);
and and17_19(wand17_19, a[17], b[19]);
and and16_19(wand16_19, a[16], b[19]);
and and15_19(wand15_19, a[15], b[19]);
and and14_19(wand14_19, a[14], b[19]);
and and13_19(wand13_19, a[13], b[19]);
and and12_19(wand12_19, a[12], b[19]);
and and11_19(wand11_19, a[11], b[19]);
and and10_19(wand10_19, a[10], b[19]);
and and9_19(wand9_19, a[9], b[19]);
and and8_19(wand8_19, a[8], b[19]);
and and7_19(wand7_19, a[7], b[19]);
and and6_19(wand6_19, a[6], b[19]);
and and5_19(wand5_19, a[5], b[19]);
and and4_19(wand4_19, a[4], b[19]);
and and3_19(wand3_19, a[3], b[19]);
and and2_19(wand2_19, a[2], b[19]);
and and1_19(wand1_19, a[1], b[19]);
and and0_19(wand0_19, a[0], b[19]);
nand nand31_20(wand31_20, a[31], b[20]);
and and30_20(wand30_20, a[30], b[20]);
and and29_20(wand29_20, a[29], b[20]);
and and28_20(wand28_20, a[28], b[20]);
and and27_20(wand27_20, a[27], b[20]);
and and26_20(wand26_20, a[26], b[20]);
and and25_20(wand25_20, a[25], b[20]);
and and24_20(wand24_20, a[24], b[20]);
and and23_20(wand23_20, a[23], b[20]);
and and22_20(wand22_20, a[22], b[20]);
and and21_20(wand21_20, a[21], b[20]);
and and20_20(wand20_20, a[20], b[20]);
and and19_20(wand19_20, a[19], b[20]);
and and18_20(wand18_20, a[18], b[20]);
and and17_20(wand17_20, a[17], b[20]);
and and16_20(wand16_20, a[16], b[20]);
and and15_20(wand15_20, a[15], b[20]);
and and14_20(wand14_20, a[14], b[20]);
and and13_20(wand13_20, a[13], b[20]);
and and12_20(wand12_20, a[12], b[20]);
and and11_20(wand11_20, a[11], b[20]);
and and10_20(wand10_20, a[10], b[20]);
and and9_20(wand9_20, a[9], b[20]);
and and8_20(wand8_20, a[8], b[20]);
and and7_20(wand7_20, a[7], b[20]);
and and6_20(wand6_20, a[6], b[20]);
and and5_20(wand5_20, a[5], b[20]);
and and4_20(wand4_20, a[4], b[20]);
and and3_20(wand3_20, a[3], b[20]);
and and2_20(wand2_20, a[2], b[20]);
and and1_20(wand1_20, a[1], b[20]);
and and0_20(wand0_20, a[0], b[20]);
nand nand31_21(wand31_21, a[31], b[21]);
and and30_21(wand30_21, a[30], b[21]);
and and29_21(wand29_21, a[29], b[21]);
and and28_21(wand28_21, a[28], b[21]);
and and27_21(wand27_21, a[27], b[21]);
and and26_21(wand26_21, a[26], b[21]);
and and25_21(wand25_21, a[25], b[21]);
and and24_21(wand24_21, a[24], b[21]);
and and23_21(wand23_21, a[23], b[21]);
and and22_21(wand22_21, a[22], b[21]);
and and21_21(wand21_21, a[21], b[21]);
and and20_21(wand20_21, a[20], b[21]);
and and19_21(wand19_21, a[19], b[21]);
and and18_21(wand18_21, a[18], b[21]);
and and17_21(wand17_21, a[17], b[21]);
and and16_21(wand16_21, a[16], b[21]);
and and15_21(wand15_21, a[15], b[21]);
and and14_21(wand14_21, a[14], b[21]);
and and13_21(wand13_21, a[13], b[21]);
and and12_21(wand12_21, a[12], b[21]);
and and11_21(wand11_21, a[11], b[21]);
and and10_21(wand10_21, a[10], b[21]);
and and9_21(wand9_21, a[9], b[21]);
and and8_21(wand8_21, a[8], b[21]);
and and7_21(wand7_21, a[7], b[21]);
and and6_21(wand6_21, a[6], b[21]);
and and5_21(wand5_21, a[5], b[21]);
and and4_21(wand4_21, a[4], b[21]);
and and3_21(wand3_21, a[3], b[21]);
and and2_21(wand2_21, a[2], b[21]);
and and1_21(wand1_21, a[1], b[21]);
and and0_21(wand0_21, a[0], b[21]);
nand nand31_22(wand31_22, a[31], b[22]);
and and30_22(wand30_22, a[30], b[22]);
and and29_22(wand29_22, a[29], b[22]);
and and28_22(wand28_22, a[28], b[22]);
and and27_22(wand27_22, a[27], b[22]);
and and26_22(wand26_22, a[26], b[22]);
and and25_22(wand25_22, a[25], b[22]);
and and24_22(wand24_22, a[24], b[22]);
and and23_22(wand23_22, a[23], b[22]);
and and22_22(wand22_22, a[22], b[22]);
and and21_22(wand21_22, a[21], b[22]);
and and20_22(wand20_22, a[20], b[22]);
and and19_22(wand19_22, a[19], b[22]);
and and18_22(wand18_22, a[18], b[22]);
and and17_22(wand17_22, a[17], b[22]);
and and16_22(wand16_22, a[16], b[22]);
and and15_22(wand15_22, a[15], b[22]);
and and14_22(wand14_22, a[14], b[22]);
and and13_22(wand13_22, a[13], b[22]);
and and12_22(wand12_22, a[12], b[22]);
and and11_22(wand11_22, a[11], b[22]);
and and10_22(wand10_22, a[10], b[22]);
and and9_22(wand9_22, a[9], b[22]);
and and8_22(wand8_22, a[8], b[22]);
and and7_22(wand7_22, a[7], b[22]);
and and6_22(wand6_22, a[6], b[22]);
and and5_22(wand5_22, a[5], b[22]);
and and4_22(wand4_22, a[4], b[22]);
and and3_22(wand3_22, a[3], b[22]);
and and2_22(wand2_22, a[2], b[22]);
and and1_22(wand1_22, a[1], b[22]);
and and0_22(wand0_22, a[0], b[22]);
nand nand31_23(wand31_23, a[31], b[23]);
and and30_23(wand30_23, a[30], b[23]);
and and29_23(wand29_23, a[29], b[23]);
and and28_23(wand28_23, a[28], b[23]);
and and27_23(wand27_23, a[27], b[23]);
and and26_23(wand26_23, a[26], b[23]);
and and25_23(wand25_23, a[25], b[23]);
and and24_23(wand24_23, a[24], b[23]);
and and23_23(wand23_23, a[23], b[23]);
and and22_23(wand22_23, a[22], b[23]);
and and21_23(wand21_23, a[21], b[23]);
and and20_23(wand20_23, a[20], b[23]);
and and19_23(wand19_23, a[19], b[23]);
and and18_23(wand18_23, a[18], b[23]);
and and17_23(wand17_23, a[17], b[23]);
and and16_23(wand16_23, a[16], b[23]);
and and15_23(wand15_23, a[15], b[23]);
and and14_23(wand14_23, a[14], b[23]);
and and13_23(wand13_23, a[13], b[23]);
and and12_23(wand12_23, a[12], b[23]);
and and11_23(wand11_23, a[11], b[23]);
and and10_23(wand10_23, a[10], b[23]);
and and9_23(wand9_23, a[9], b[23]);
and and8_23(wand8_23, a[8], b[23]);
and and7_23(wand7_23, a[7], b[23]);
and and6_23(wand6_23, a[6], b[23]);
and and5_23(wand5_23, a[5], b[23]);
and and4_23(wand4_23, a[4], b[23]);
and and3_23(wand3_23, a[3], b[23]);
and and2_23(wand2_23, a[2], b[23]);
and and1_23(wand1_23, a[1], b[23]);
and and0_23(wand0_23, a[0], b[23]);
nand nand31_24(wand31_24, a[31], b[24]);
and and30_24(wand30_24, a[30], b[24]);
and and29_24(wand29_24, a[29], b[24]);
and and28_24(wand28_24, a[28], b[24]);
and and27_24(wand27_24, a[27], b[24]);
and and26_24(wand26_24, a[26], b[24]);
and and25_24(wand25_24, a[25], b[24]);
and and24_24(wand24_24, a[24], b[24]);
and and23_24(wand23_24, a[23], b[24]);
and and22_24(wand22_24, a[22], b[24]);
and and21_24(wand21_24, a[21], b[24]);
and and20_24(wand20_24, a[20], b[24]);
and and19_24(wand19_24, a[19], b[24]);
and and18_24(wand18_24, a[18], b[24]);
and and17_24(wand17_24, a[17], b[24]);
and and16_24(wand16_24, a[16], b[24]);
and and15_24(wand15_24, a[15], b[24]);
and and14_24(wand14_24, a[14], b[24]);
and and13_24(wand13_24, a[13], b[24]);
and and12_24(wand12_24, a[12], b[24]);
and and11_24(wand11_24, a[11], b[24]);
and and10_24(wand10_24, a[10], b[24]);
and and9_24(wand9_24, a[9], b[24]);
and and8_24(wand8_24, a[8], b[24]);
and and7_24(wand7_24, a[7], b[24]);
and and6_24(wand6_24, a[6], b[24]);
and and5_24(wand5_24, a[5], b[24]);
and and4_24(wand4_24, a[4], b[24]);
and and3_24(wand3_24, a[3], b[24]);
and and2_24(wand2_24, a[2], b[24]);
and and1_24(wand1_24, a[1], b[24]);
and and0_24(wand0_24, a[0], b[24]);
nand nand31_25(wand31_25, a[31], b[25]);
and and30_25(wand30_25, a[30], b[25]);
and and29_25(wand29_25, a[29], b[25]);
and and28_25(wand28_25, a[28], b[25]);
and and27_25(wand27_25, a[27], b[25]);
and and26_25(wand26_25, a[26], b[25]);
and and25_25(wand25_25, a[25], b[25]);
and and24_25(wand24_25, a[24], b[25]);
and and23_25(wand23_25, a[23], b[25]);
and and22_25(wand22_25, a[22], b[25]);
and and21_25(wand21_25, a[21], b[25]);
and and20_25(wand20_25, a[20], b[25]);
and and19_25(wand19_25, a[19], b[25]);
and and18_25(wand18_25, a[18], b[25]);
and and17_25(wand17_25, a[17], b[25]);
and and16_25(wand16_25, a[16], b[25]);
and and15_25(wand15_25, a[15], b[25]);
and and14_25(wand14_25, a[14], b[25]);
and and13_25(wand13_25, a[13], b[25]);
and and12_25(wand12_25, a[12], b[25]);
and and11_25(wand11_25, a[11], b[25]);
and and10_25(wand10_25, a[10], b[25]);
and and9_25(wand9_25, a[9], b[25]);
and and8_25(wand8_25, a[8], b[25]);
and and7_25(wand7_25, a[7], b[25]);
and and6_25(wand6_25, a[6], b[25]);
and and5_25(wand5_25, a[5], b[25]);
and and4_25(wand4_25, a[4], b[25]);
and and3_25(wand3_25, a[3], b[25]);
and and2_25(wand2_25, a[2], b[25]);
and and1_25(wand1_25, a[1], b[25]);
and and0_25(wand0_25, a[0], b[25]);
nand nand31_26(wand31_26, a[31], b[26]);
and and30_26(wand30_26, a[30], b[26]);
and and29_26(wand29_26, a[29], b[26]);
and and28_26(wand28_26, a[28], b[26]);
and and27_26(wand27_26, a[27], b[26]);
and and26_26(wand26_26, a[26], b[26]);
and and25_26(wand25_26, a[25], b[26]);
and and24_26(wand24_26, a[24], b[26]);
and and23_26(wand23_26, a[23], b[26]);
and and22_26(wand22_26, a[22], b[26]);
and and21_26(wand21_26, a[21], b[26]);
and and20_26(wand20_26, a[20], b[26]);
and and19_26(wand19_26, a[19], b[26]);
and and18_26(wand18_26, a[18], b[26]);
and and17_26(wand17_26, a[17], b[26]);
and and16_26(wand16_26, a[16], b[26]);
and and15_26(wand15_26, a[15], b[26]);
and and14_26(wand14_26, a[14], b[26]);
and and13_26(wand13_26, a[13], b[26]);
and and12_26(wand12_26, a[12], b[26]);
and and11_26(wand11_26, a[11], b[26]);
and and10_26(wand10_26, a[10], b[26]);
and and9_26(wand9_26, a[9], b[26]);
and and8_26(wand8_26, a[8], b[26]);
and and7_26(wand7_26, a[7], b[26]);
and and6_26(wand6_26, a[6], b[26]);
and and5_26(wand5_26, a[5], b[26]);
and and4_26(wand4_26, a[4], b[26]);
and and3_26(wand3_26, a[3], b[26]);
and and2_26(wand2_26, a[2], b[26]);
and and1_26(wand1_26, a[1], b[26]);
and and0_26(wand0_26, a[0], b[26]);
nand nand31_27(wand31_27, a[31], b[27]);
and and30_27(wand30_27, a[30], b[27]);
and and29_27(wand29_27, a[29], b[27]);
and and28_27(wand28_27, a[28], b[27]);
and and27_27(wand27_27, a[27], b[27]);
and and26_27(wand26_27, a[26], b[27]);
and and25_27(wand25_27, a[25], b[27]);
and and24_27(wand24_27, a[24], b[27]);
and and23_27(wand23_27, a[23], b[27]);
and and22_27(wand22_27, a[22], b[27]);
and and21_27(wand21_27, a[21], b[27]);
and and20_27(wand20_27, a[20], b[27]);
and and19_27(wand19_27, a[19], b[27]);
and and18_27(wand18_27, a[18], b[27]);
and and17_27(wand17_27, a[17], b[27]);
and and16_27(wand16_27, a[16], b[27]);
and and15_27(wand15_27, a[15], b[27]);
and and14_27(wand14_27, a[14], b[27]);
and and13_27(wand13_27, a[13], b[27]);
and and12_27(wand12_27, a[12], b[27]);
and and11_27(wand11_27, a[11], b[27]);
and and10_27(wand10_27, a[10], b[27]);
and and9_27(wand9_27, a[9], b[27]);
and and8_27(wand8_27, a[8], b[27]);
and and7_27(wand7_27, a[7], b[27]);
and and6_27(wand6_27, a[6], b[27]);
and and5_27(wand5_27, a[5], b[27]);
and and4_27(wand4_27, a[4], b[27]);
and and3_27(wand3_27, a[3], b[27]);
and and2_27(wand2_27, a[2], b[27]);
and and1_27(wand1_27, a[1], b[27]);
and and0_27(wand0_27, a[0], b[27]);
nand nand31_28(wand31_28, a[31], b[28]);
and and30_28(wand30_28, a[30], b[28]);
and and29_28(wand29_28, a[29], b[28]);
and and28_28(wand28_28, a[28], b[28]);
and and27_28(wand27_28, a[27], b[28]);
and and26_28(wand26_28, a[26], b[28]);
and and25_28(wand25_28, a[25], b[28]);
and and24_28(wand24_28, a[24], b[28]);
and and23_28(wand23_28, a[23], b[28]);
and and22_28(wand22_28, a[22], b[28]);
and and21_28(wand21_28, a[21], b[28]);
and and20_28(wand20_28, a[20], b[28]);
and and19_28(wand19_28, a[19], b[28]);
and and18_28(wand18_28, a[18], b[28]);
and and17_28(wand17_28, a[17], b[28]);
and and16_28(wand16_28, a[16], b[28]);
and and15_28(wand15_28, a[15], b[28]);
and and14_28(wand14_28, a[14], b[28]);
and and13_28(wand13_28, a[13], b[28]);
and and12_28(wand12_28, a[12], b[28]);
and and11_28(wand11_28, a[11], b[28]);
and and10_28(wand10_28, a[10], b[28]);
and and9_28(wand9_28, a[9], b[28]);
and and8_28(wand8_28, a[8], b[28]);
and and7_28(wand7_28, a[7], b[28]);
and and6_28(wand6_28, a[6], b[28]);
and and5_28(wand5_28, a[5], b[28]);
and and4_28(wand4_28, a[4], b[28]);
and and3_28(wand3_28, a[3], b[28]);
and and2_28(wand2_28, a[2], b[28]);
and and1_28(wand1_28, a[1], b[28]);
and and0_28(wand0_28, a[0], b[28]);
nand nand31_29(wand31_29, a[31], b[29]);
and and30_29(wand30_29, a[30], b[29]);
and and29_29(wand29_29, a[29], b[29]);
and and28_29(wand28_29, a[28], b[29]);
and and27_29(wand27_29, a[27], b[29]);
and and26_29(wand26_29, a[26], b[29]);
and and25_29(wand25_29, a[25], b[29]);
and and24_29(wand24_29, a[24], b[29]);
and and23_29(wand23_29, a[23], b[29]);
and and22_29(wand22_29, a[22], b[29]);
and and21_29(wand21_29, a[21], b[29]);
and and20_29(wand20_29, a[20], b[29]);
and and19_29(wand19_29, a[19], b[29]);
and and18_29(wand18_29, a[18], b[29]);
and and17_29(wand17_29, a[17], b[29]);
and and16_29(wand16_29, a[16], b[29]);
and and15_29(wand15_29, a[15], b[29]);
and and14_29(wand14_29, a[14], b[29]);
and and13_29(wand13_29, a[13], b[29]);
and and12_29(wand12_29, a[12], b[29]);
and and11_29(wand11_29, a[11], b[29]);
and and10_29(wand10_29, a[10], b[29]);
and and9_29(wand9_29, a[9], b[29]);
and and8_29(wand8_29, a[8], b[29]);
and and7_29(wand7_29, a[7], b[29]);
and and6_29(wand6_29, a[6], b[29]);
and and5_29(wand5_29, a[5], b[29]);
and and4_29(wand4_29, a[4], b[29]);
and and3_29(wand3_29, a[3], b[29]);
and and2_29(wand2_29, a[2], b[29]);
and and1_29(wand1_29, a[1], b[29]);
and and0_29(wand0_29, a[0], b[29]);
nand nand31_30(wand31_30, a[31], b[30]);
and and30_30(wand30_30, a[30], b[30]);
and and29_30(wand29_30, a[29], b[30]);
and and28_30(wand28_30, a[28], b[30]);
and and27_30(wand27_30, a[27], b[30]);
and and26_30(wand26_30, a[26], b[30]);
and and25_30(wand25_30, a[25], b[30]);
and and24_30(wand24_30, a[24], b[30]);
and and23_30(wand23_30, a[23], b[30]);
and and22_30(wand22_30, a[22], b[30]);
and and21_30(wand21_30, a[21], b[30]);
and and20_30(wand20_30, a[20], b[30]);
and and19_30(wand19_30, a[19], b[30]);
and and18_30(wand18_30, a[18], b[30]);
and and17_30(wand17_30, a[17], b[30]);
and and16_30(wand16_30, a[16], b[30]);
and and15_30(wand15_30, a[15], b[30]);
and and14_30(wand14_30, a[14], b[30]);
and and13_30(wand13_30, a[13], b[30]);
and and12_30(wand12_30, a[12], b[30]);
and and11_30(wand11_30, a[11], b[30]);
and and10_30(wand10_30, a[10], b[30]);
and and9_30(wand9_30, a[9], b[30]);
and and8_30(wand8_30, a[8], b[30]);
and and7_30(wand7_30, a[7], b[30]);
and and6_30(wand6_30, a[6], b[30]);
and and5_30(wand5_30, a[5], b[30]);
and and4_30(wand4_30, a[4], b[30]);
and and3_30(wand3_30, a[3], b[30]);
and and2_30(wand2_30, a[2], b[30]);
and and1_30(wand1_30, a[1], b[30]);
and and0_30(wand0_30, a[0], b[30]);
and and31_31(wand31_31, a[31], b[31]);
nand nand30_31(wand30_31, a[30], b[31]);
nand nand29_31(wand29_31, a[29], b[31]);
nand nand28_31(wand28_31, a[28], b[31]);
nand nand27_31(wand27_31, a[27], b[31]);
nand nand26_31(wand26_31, a[26], b[31]);
nand nand25_31(wand25_31, a[25], b[31]);
nand nand24_31(wand24_31, a[24], b[31]);
nand nand23_31(wand23_31, a[23], b[31]);
nand nand22_31(wand22_31, a[22], b[31]);
nand nand21_31(wand21_31, a[21], b[31]);
nand nand20_31(wand20_31, a[20], b[31]);
nand nand19_31(wand19_31, a[19], b[31]);
nand nand18_31(wand18_31, a[18], b[31]);
nand nand17_31(wand17_31, a[17], b[31]);
nand nand16_31(wand16_31, a[16], b[31]);
nand nand15_31(wand15_31, a[15], b[31]);
nand nand14_31(wand14_31, a[14], b[31]);
nand nand13_31(wand13_31, a[13], b[31]);
nand nand12_31(wand12_31, a[12], b[31]);
nand nand11_31(wand11_31, a[11], b[31]);
nand nand10_31(wand10_31, a[10], b[31]);
nand nand9_31(wand9_31, a[9], b[31]);
nand nand8_31(wand8_31, a[8], b[31]);
nand nand7_31(wand7_31, a[7], b[31]);
nand nand6_31(wand6_31, a[6], b[31]);
nand nand5_31(wand5_31, a[5], b[31]);
nand nand4_31(wand4_31, a[4], b[31]);
nand nand3_31(wand3_31, a[3], b[31]);
nand nand2_31(wand2_31, a[2], b[31]);
nand nand1_31(wand1_31, a[1], b[31]);
nand nand0_31(wand0_31, a[0], b[31]);


assign ws0b0n0_30 = wand31_2;
adder_full fa0(.sum(ws0b0n0_31), .c_out(ws0b0n1_30), .a(wand31_1), .b(wand30_2), .c_in(1'b1));
adder_full fa1(.sum(ws0b0n0_32), .c_out(ws0b0n1_31), .a(wand31_0), .b(wand30_1), .c_in(wand29_2));
adder_full fa2(.sum(ws0b0n0_33), .c_out(ws0b0n1_32), .a(wand30_0), .b(wand29_1), .c_in(wand28_2));
adder_full fa3(.sum(ws0b0n0_34), .c_out(ws0b0n1_33), .a(wand29_0), .b(wand28_1), .c_in(wand27_2));
adder_full fa4(.sum(ws0b0n0_35), .c_out(ws0b0n1_34), .a(wand28_0), .b(wand27_1), .c_in(wand26_2));
adder_full fa5(.sum(ws0b0n0_36), .c_out(ws0b0n1_35), .a(wand27_0), .b(wand26_1), .c_in(wand25_2));
adder_full fa6(.sum(ws0b0n0_37), .c_out(ws0b0n1_36), .a(wand26_0), .b(wand25_1), .c_in(wand24_2));
adder_full fa7(.sum(ws0b0n0_38), .c_out(ws0b0n1_37), .a(wand25_0), .b(wand24_1), .c_in(wand23_2));
adder_full fa8(.sum(ws0b0n0_39), .c_out(ws0b0n1_38), .a(wand24_0), .b(wand23_1), .c_in(wand22_2));
adder_full fa9(.sum(ws0b0n0_40), .c_out(ws0b0n1_39), .a(wand23_0), .b(wand22_1), .c_in(wand21_2));
adder_full fa10(.sum(ws0b0n0_41), .c_out(ws0b0n1_40), .a(wand22_0), .b(wand21_1), .c_in(wand20_2));
adder_full fa11(.sum(ws0b0n0_42), .c_out(ws0b0n1_41), .a(wand21_0), .b(wand20_1), .c_in(wand19_2));
adder_full fa12(.sum(ws0b0n0_43), .c_out(ws0b0n1_42), .a(wand20_0), .b(wand19_1), .c_in(wand18_2));
adder_full fa13(.sum(ws0b0n0_44), .c_out(ws0b0n1_43), .a(wand19_0), .b(wand18_1), .c_in(wand17_2));
adder_full fa14(.sum(ws0b0n0_45), .c_out(ws0b0n1_44), .a(wand18_0), .b(wand17_1), .c_in(wand16_2));
adder_full fa15(.sum(ws0b0n0_46), .c_out(ws0b0n1_45), .a(wand17_0), .b(wand16_1), .c_in(wand15_2));
adder_full fa16(.sum(ws0b0n0_47), .c_out(ws0b0n1_46), .a(wand16_0), .b(wand15_1), .c_in(wand14_2));
adder_full fa17(.sum(ws0b0n0_48), .c_out(ws0b0n1_47), .a(wand15_0), .b(wand14_1), .c_in(wand13_2));
adder_full fa18(.sum(ws0b0n0_49), .c_out(ws0b0n1_48), .a(wand14_0), .b(wand13_1), .c_in(wand12_2));
adder_full fa19(.sum(ws0b0n0_50), .c_out(ws0b0n1_49), .a(wand13_0), .b(wand12_1), .c_in(wand11_2));
adder_full fa20(.sum(ws0b0n0_51), .c_out(ws0b0n1_50), .a(wand12_0), .b(wand11_1), .c_in(wand10_2));
adder_full fa21(.sum(ws0b0n0_52), .c_out(ws0b0n1_51), .a(wand11_0), .b(wand10_1), .c_in(wand9_2));
adder_full fa22(.sum(ws0b0n0_53), .c_out(ws0b0n1_52), .a(wand10_0), .b(wand9_1), .c_in(wand8_2));
adder_full fa23(.sum(ws0b0n0_54), .c_out(ws0b0n1_53), .a(wand9_0), .b(wand8_1), .c_in(wand7_2));
adder_full fa24(.sum(ws0b0n0_55), .c_out(ws0b0n1_54), .a(wand8_0), .b(wand7_1), .c_in(wand6_2));
adder_full fa25(.sum(ws0b0n0_56), .c_out(ws0b0n1_55), .a(wand7_0), .b(wand6_1), .c_in(wand5_2));
adder_full fa26(.sum(ws0b0n0_57), .c_out(ws0b0n1_56), .a(wand6_0), .b(wand5_1), .c_in(wand4_2));
adder_full fa27(.sum(ws0b0n0_58), .c_out(ws0b0n1_57), .a(wand5_0), .b(wand4_1), .c_in(wand3_2));
adder_full fa28(.sum(ws0b0n0_59), .c_out(ws0b0n1_58), .a(wand4_0), .b(wand3_1), .c_in(wand2_2));
adder_full fa29(.sum(ws0b0n0_60), .c_out(ws0b0n1_59), .a(wand3_0), .b(wand2_1), .c_in(wand1_2));
adder_full fa30(.sum(ws0b0n0_61), .c_out(ws0b0n1_60), .a(wand2_0), .b(wand1_1), .c_in(wand0_2));
adder_half ha0(.sum(ws0b0n0_62), .c_out(ws0b0n1_61), .a(wand1_0), .b(wand0_1));
assign ws0b0n0_63 = wand0_0;
assign ws0b1n0_27 = wand31_5;
adder_half ha1(.sum(ws0b1n0_28), .c_out(ws0b1n1_27), .a(wand31_4), .b(wand30_5));
adder_full fa31(.sum(ws0b1n0_29), .c_out(ws0b1n1_28), .a(wand31_3), .b(wand30_4), .c_in(wand29_5));
adder_full fa32(.sum(ws0b1n0_30), .c_out(ws0b1n1_29), .a(wand30_3), .b(wand29_4), .c_in(wand28_5));
adder_full fa33(.sum(ws0b1n0_31), .c_out(ws0b1n1_30), .a(wand29_3), .b(wand28_4), .c_in(wand27_5));
adder_full fa34(.sum(ws0b1n0_32), .c_out(ws0b1n1_31), .a(wand28_3), .b(wand27_4), .c_in(wand26_5));
adder_full fa35(.sum(ws0b1n0_33), .c_out(ws0b1n1_32), .a(wand27_3), .b(wand26_4), .c_in(wand25_5));
adder_full fa36(.sum(ws0b1n0_34), .c_out(ws0b1n1_33), .a(wand26_3), .b(wand25_4), .c_in(wand24_5));
adder_full fa37(.sum(ws0b1n0_35), .c_out(ws0b1n1_34), .a(wand25_3), .b(wand24_4), .c_in(wand23_5));
adder_full fa38(.sum(ws0b1n0_36), .c_out(ws0b1n1_35), .a(wand24_3), .b(wand23_4), .c_in(wand22_5));
adder_full fa39(.sum(ws0b1n0_37), .c_out(ws0b1n1_36), .a(wand23_3), .b(wand22_4), .c_in(wand21_5));
adder_full fa40(.sum(ws0b1n0_38), .c_out(ws0b1n1_37), .a(wand22_3), .b(wand21_4), .c_in(wand20_5));
adder_full fa41(.sum(ws0b1n0_39), .c_out(ws0b1n1_38), .a(wand21_3), .b(wand20_4), .c_in(wand19_5));
adder_full fa42(.sum(ws0b1n0_40), .c_out(ws0b1n1_39), .a(wand20_3), .b(wand19_4), .c_in(wand18_5));
adder_full fa43(.sum(ws0b1n0_41), .c_out(ws0b1n1_40), .a(wand19_3), .b(wand18_4), .c_in(wand17_5));
adder_full fa44(.sum(ws0b1n0_42), .c_out(ws0b1n1_41), .a(wand18_3), .b(wand17_4), .c_in(wand16_5));
adder_full fa45(.sum(ws0b1n0_43), .c_out(ws0b1n1_42), .a(wand17_3), .b(wand16_4), .c_in(wand15_5));
adder_full fa46(.sum(ws0b1n0_44), .c_out(ws0b1n1_43), .a(wand16_3), .b(wand15_4), .c_in(wand14_5));
adder_full fa47(.sum(ws0b1n0_45), .c_out(ws0b1n1_44), .a(wand15_3), .b(wand14_4), .c_in(wand13_5));
adder_full fa48(.sum(ws0b1n0_46), .c_out(ws0b1n1_45), .a(wand14_3), .b(wand13_4), .c_in(wand12_5));
adder_full fa49(.sum(ws0b1n0_47), .c_out(ws0b1n1_46), .a(wand13_3), .b(wand12_4), .c_in(wand11_5));
adder_full fa50(.sum(ws0b1n0_48), .c_out(ws0b1n1_47), .a(wand12_3), .b(wand11_4), .c_in(wand10_5));
adder_full fa51(.sum(ws0b1n0_49), .c_out(ws0b1n1_48), .a(wand11_3), .b(wand10_4), .c_in(wand9_5));
adder_full fa52(.sum(ws0b1n0_50), .c_out(ws0b1n1_49), .a(wand10_3), .b(wand9_4), .c_in(wand8_5));
adder_full fa53(.sum(ws0b1n0_51), .c_out(ws0b1n1_50), .a(wand9_3), .b(wand8_4), .c_in(wand7_5));
adder_full fa54(.sum(ws0b1n0_52), .c_out(ws0b1n1_51), .a(wand8_3), .b(wand7_4), .c_in(wand6_5));
adder_full fa55(.sum(ws0b1n0_53), .c_out(ws0b1n1_52), .a(wand7_3), .b(wand6_4), .c_in(wand5_5));
adder_full fa56(.sum(ws0b1n0_54), .c_out(ws0b1n1_53), .a(wand6_3), .b(wand5_4), .c_in(wand4_5));
adder_full fa57(.sum(ws0b1n0_55), .c_out(ws0b1n1_54), .a(wand5_3), .b(wand4_4), .c_in(wand3_5));
adder_full fa58(.sum(ws0b1n0_56), .c_out(ws0b1n1_55), .a(wand4_3), .b(wand3_4), .c_in(wand2_5));
adder_full fa59(.sum(ws0b1n0_57), .c_out(ws0b1n1_56), .a(wand3_3), .b(wand2_4), .c_in(wand1_5));
adder_full fa60(.sum(ws0b1n0_58), .c_out(ws0b1n1_57), .a(wand2_3), .b(wand1_4), .c_in(wand0_5));
adder_half ha2(.sum(ws0b1n0_59), .c_out(ws0b1n1_58), .a(wand1_3), .b(wand0_4));
assign ws0b1n0_60 = wand0_3;
assign ws0b2n0_24 = wand31_8;
adder_half ha3(.sum(ws0b2n0_25), .c_out(ws0b2n1_24), .a(wand31_7), .b(wand30_8));
adder_full fa61(.sum(ws0b2n0_26), .c_out(ws0b2n1_25), .a(wand31_6), .b(wand30_7), .c_in(wand29_8));
adder_full fa62(.sum(ws0b2n0_27), .c_out(ws0b2n1_26), .a(wand30_6), .b(wand29_7), .c_in(wand28_8));
adder_full fa63(.sum(ws0b2n0_28), .c_out(ws0b2n1_27), .a(wand29_6), .b(wand28_7), .c_in(wand27_8));
adder_full fa64(.sum(ws0b2n0_29), .c_out(ws0b2n1_28), .a(wand28_6), .b(wand27_7), .c_in(wand26_8));
adder_full fa65(.sum(ws0b2n0_30), .c_out(ws0b2n1_29), .a(wand27_6), .b(wand26_7), .c_in(wand25_8));
adder_full fa66(.sum(ws0b2n0_31), .c_out(ws0b2n1_30), .a(wand26_6), .b(wand25_7), .c_in(wand24_8));
adder_full fa67(.sum(ws0b2n0_32), .c_out(ws0b2n1_31), .a(wand25_6), .b(wand24_7), .c_in(wand23_8));
adder_full fa68(.sum(ws0b2n0_33), .c_out(ws0b2n1_32), .a(wand24_6), .b(wand23_7), .c_in(wand22_8));
adder_full fa69(.sum(ws0b2n0_34), .c_out(ws0b2n1_33), .a(wand23_6), .b(wand22_7), .c_in(wand21_8));
adder_full fa70(.sum(ws0b2n0_35), .c_out(ws0b2n1_34), .a(wand22_6), .b(wand21_7), .c_in(wand20_8));
adder_full fa71(.sum(ws0b2n0_36), .c_out(ws0b2n1_35), .a(wand21_6), .b(wand20_7), .c_in(wand19_8));
adder_full fa72(.sum(ws0b2n0_37), .c_out(ws0b2n1_36), .a(wand20_6), .b(wand19_7), .c_in(wand18_8));
adder_full fa73(.sum(ws0b2n0_38), .c_out(ws0b2n1_37), .a(wand19_6), .b(wand18_7), .c_in(wand17_8));
adder_full fa74(.sum(ws0b2n0_39), .c_out(ws0b2n1_38), .a(wand18_6), .b(wand17_7), .c_in(wand16_8));
adder_full fa75(.sum(ws0b2n0_40), .c_out(ws0b2n1_39), .a(wand17_6), .b(wand16_7), .c_in(wand15_8));
adder_full fa76(.sum(ws0b2n0_41), .c_out(ws0b2n1_40), .a(wand16_6), .b(wand15_7), .c_in(wand14_8));
adder_full fa77(.sum(ws0b2n0_42), .c_out(ws0b2n1_41), .a(wand15_6), .b(wand14_7), .c_in(wand13_8));
adder_full fa78(.sum(ws0b2n0_43), .c_out(ws0b2n1_42), .a(wand14_6), .b(wand13_7), .c_in(wand12_8));
adder_full fa79(.sum(ws0b2n0_44), .c_out(ws0b2n1_43), .a(wand13_6), .b(wand12_7), .c_in(wand11_8));
adder_full fa80(.sum(ws0b2n0_45), .c_out(ws0b2n1_44), .a(wand12_6), .b(wand11_7), .c_in(wand10_8));
adder_full fa81(.sum(ws0b2n0_46), .c_out(ws0b2n1_45), .a(wand11_6), .b(wand10_7), .c_in(wand9_8));
adder_full fa82(.sum(ws0b2n0_47), .c_out(ws0b2n1_46), .a(wand10_6), .b(wand9_7), .c_in(wand8_8));
adder_full fa83(.sum(ws0b2n0_48), .c_out(ws0b2n1_47), .a(wand9_6), .b(wand8_7), .c_in(wand7_8));
adder_full fa84(.sum(ws0b2n0_49), .c_out(ws0b2n1_48), .a(wand8_6), .b(wand7_7), .c_in(wand6_8));
adder_full fa85(.sum(ws0b2n0_50), .c_out(ws0b2n1_49), .a(wand7_6), .b(wand6_7), .c_in(wand5_8));
adder_full fa86(.sum(ws0b2n0_51), .c_out(ws0b2n1_50), .a(wand6_6), .b(wand5_7), .c_in(wand4_8));
adder_full fa87(.sum(ws0b2n0_52), .c_out(ws0b2n1_51), .a(wand5_6), .b(wand4_7), .c_in(wand3_8));
adder_full fa88(.sum(ws0b2n0_53), .c_out(ws0b2n1_52), .a(wand4_6), .b(wand3_7), .c_in(wand2_8));
adder_full fa89(.sum(ws0b2n0_54), .c_out(ws0b2n1_53), .a(wand3_6), .b(wand2_7), .c_in(wand1_8));
adder_full fa90(.sum(ws0b2n0_55), .c_out(ws0b2n1_54), .a(wand2_6), .b(wand1_7), .c_in(wand0_8));
adder_half ha4(.sum(ws0b2n0_56), .c_out(ws0b2n1_55), .a(wand1_6), .b(wand0_7));
assign ws0b2n0_57 = wand0_6;
assign ws0b3n0_21 = wand31_11;
adder_half ha5(.sum(ws0b3n0_22), .c_out(ws0b3n1_21), .a(wand31_10), .b(wand30_11));
adder_full fa91(.sum(ws0b3n0_23), .c_out(ws0b3n1_22), .a(wand31_9), .b(wand30_10), .c_in(wand29_11));
adder_full fa92(.sum(ws0b3n0_24), .c_out(ws0b3n1_23), .a(wand30_9), .b(wand29_10), .c_in(wand28_11));
adder_full fa93(.sum(ws0b3n0_25), .c_out(ws0b3n1_24), .a(wand29_9), .b(wand28_10), .c_in(wand27_11));
adder_full fa94(.sum(ws0b3n0_26), .c_out(ws0b3n1_25), .a(wand28_9), .b(wand27_10), .c_in(wand26_11));
adder_full fa95(.sum(ws0b3n0_27), .c_out(ws0b3n1_26), .a(wand27_9), .b(wand26_10), .c_in(wand25_11));
adder_full fa96(.sum(ws0b3n0_28), .c_out(ws0b3n1_27), .a(wand26_9), .b(wand25_10), .c_in(wand24_11));
adder_full fa97(.sum(ws0b3n0_29), .c_out(ws0b3n1_28), .a(wand25_9), .b(wand24_10), .c_in(wand23_11));
adder_full fa98(.sum(ws0b3n0_30), .c_out(ws0b3n1_29), .a(wand24_9), .b(wand23_10), .c_in(wand22_11));
adder_full fa99(.sum(ws0b3n0_31), .c_out(ws0b3n1_30), .a(wand23_9), .b(wand22_10), .c_in(wand21_11));
adder_full fa100(.sum(ws0b3n0_32), .c_out(ws0b3n1_31), .a(wand22_9), .b(wand21_10), .c_in(wand20_11));
adder_full fa101(.sum(ws0b3n0_33), .c_out(ws0b3n1_32), .a(wand21_9), .b(wand20_10), .c_in(wand19_11));
adder_full fa102(.sum(ws0b3n0_34), .c_out(ws0b3n1_33), .a(wand20_9), .b(wand19_10), .c_in(wand18_11));
adder_full fa103(.sum(ws0b3n0_35), .c_out(ws0b3n1_34), .a(wand19_9), .b(wand18_10), .c_in(wand17_11));
adder_full fa104(.sum(ws0b3n0_36), .c_out(ws0b3n1_35), .a(wand18_9), .b(wand17_10), .c_in(wand16_11));
adder_full fa105(.sum(ws0b3n0_37), .c_out(ws0b3n1_36), .a(wand17_9), .b(wand16_10), .c_in(wand15_11));
adder_full fa106(.sum(ws0b3n0_38), .c_out(ws0b3n1_37), .a(wand16_9), .b(wand15_10), .c_in(wand14_11));
adder_full fa107(.sum(ws0b3n0_39), .c_out(ws0b3n1_38), .a(wand15_9), .b(wand14_10), .c_in(wand13_11));
adder_full fa108(.sum(ws0b3n0_40), .c_out(ws0b3n1_39), .a(wand14_9), .b(wand13_10), .c_in(wand12_11));
adder_full fa109(.sum(ws0b3n0_41), .c_out(ws0b3n1_40), .a(wand13_9), .b(wand12_10), .c_in(wand11_11));
adder_full fa110(.sum(ws0b3n0_42), .c_out(ws0b3n1_41), .a(wand12_9), .b(wand11_10), .c_in(wand10_11));
adder_full fa111(.sum(ws0b3n0_43), .c_out(ws0b3n1_42), .a(wand11_9), .b(wand10_10), .c_in(wand9_11));
adder_full fa112(.sum(ws0b3n0_44), .c_out(ws0b3n1_43), .a(wand10_9), .b(wand9_10), .c_in(wand8_11));
adder_full fa113(.sum(ws0b3n0_45), .c_out(ws0b3n1_44), .a(wand9_9), .b(wand8_10), .c_in(wand7_11));
adder_full fa114(.sum(ws0b3n0_46), .c_out(ws0b3n1_45), .a(wand8_9), .b(wand7_10), .c_in(wand6_11));
adder_full fa115(.sum(ws0b3n0_47), .c_out(ws0b3n1_46), .a(wand7_9), .b(wand6_10), .c_in(wand5_11));
adder_full fa116(.sum(ws0b3n0_48), .c_out(ws0b3n1_47), .a(wand6_9), .b(wand5_10), .c_in(wand4_11));
adder_full fa117(.sum(ws0b3n0_49), .c_out(ws0b3n1_48), .a(wand5_9), .b(wand4_10), .c_in(wand3_11));
adder_full fa118(.sum(ws0b3n0_50), .c_out(ws0b3n1_49), .a(wand4_9), .b(wand3_10), .c_in(wand2_11));
adder_full fa119(.sum(ws0b3n0_51), .c_out(ws0b3n1_50), .a(wand3_9), .b(wand2_10), .c_in(wand1_11));
adder_full fa120(.sum(ws0b3n0_52), .c_out(ws0b3n1_51), .a(wand2_9), .b(wand1_10), .c_in(wand0_11));
adder_half ha6(.sum(ws0b3n0_53), .c_out(ws0b3n1_52), .a(wand1_9), .b(wand0_10));
assign ws0b3n0_54 = wand0_9;
assign ws0b4n0_18 = wand31_14;
adder_half ha7(.sum(ws0b4n0_19), .c_out(ws0b4n1_18), .a(wand31_13), .b(wand30_14));
adder_full fa121(.sum(ws0b4n0_20), .c_out(ws0b4n1_19), .a(wand31_12), .b(wand30_13), .c_in(wand29_14));
adder_full fa122(.sum(ws0b4n0_21), .c_out(ws0b4n1_20), .a(wand30_12), .b(wand29_13), .c_in(wand28_14));
adder_full fa123(.sum(ws0b4n0_22), .c_out(ws0b4n1_21), .a(wand29_12), .b(wand28_13), .c_in(wand27_14));
adder_full fa124(.sum(ws0b4n0_23), .c_out(ws0b4n1_22), .a(wand28_12), .b(wand27_13), .c_in(wand26_14));
adder_full fa125(.sum(ws0b4n0_24), .c_out(ws0b4n1_23), .a(wand27_12), .b(wand26_13), .c_in(wand25_14));
adder_full fa126(.sum(ws0b4n0_25), .c_out(ws0b4n1_24), .a(wand26_12), .b(wand25_13), .c_in(wand24_14));
adder_full fa127(.sum(ws0b4n0_26), .c_out(ws0b4n1_25), .a(wand25_12), .b(wand24_13), .c_in(wand23_14));
adder_full fa128(.sum(ws0b4n0_27), .c_out(ws0b4n1_26), .a(wand24_12), .b(wand23_13), .c_in(wand22_14));
adder_full fa129(.sum(ws0b4n0_28), .c_out(ws0b4n1_27), .a(wand23_12), .b(wand22_13), .c_in(wand21_14));
adder_full fa130(.sum(ws0b4n0_29), .c_out(ws0b4n1_28), .a(wand22_12), .b(wand21_13), .c_in(wand20_14));
adder_full fa131(.sum(ws0b4n0_30), .c_out(ws0b4n1_29), .a(wand21_12), .b(wand20_13), .c_in(wand19_14));
adder_full fa132(.sum(ws0b4n0_31), .c_out(ws0b4n1_30), .a(wand20_12), .b(wand19_13), .c_in(wand18_14));
adder_full fa133(.sum(ws0b4n0_32), .c_out(ws0b4n1_31), .a(wand19_12), .b(wand18_13), .c_in(wand17_14));
adder_full fa134(.sum(ws0b4n0_33), .c_out(ws0b4n1_32), .a(wand18_12), .b(wand17_13), .c_in(wand16_14));
adder_full fa135(.sum(ws0b4n0_34), .c_out(ws0b4n1_33), .a(wand17_12), .b(wand16_13), .c_in(wand15_14));
adder_full fa136(.sum(ws0b4n0_35), .c_out(ws0b4n1_34), .a(wand16_12), .b(wand15_13), .c_in(wand14_14));
adder_full fa137(.sum(ws0b4n0_36), .c_out(ws0b4n1_35), .a(wand15_12), .b(wand14_13), .c_in(wand13_14));
adder_full fa138(.sum(ws0b4n0_37), .c_out(ws0b4n1_36), .a(wand14_12), .b(wand13_13), .c_in(wand12_14));
adder_full fa139(.sum(ws0b4n0_38), .c_out(ws0b4n1_37), .a(wand13_12), .b(wand12_13), .c_in(wand11_14));
adder_full fa140(.sum(ws0b4n0_39), .c_out(ws0b4n1_38), .a(wand12_12), .b(wand11_13), .c_in(wand10_14));
adder_full fa141(.sum(ws0b4n0_40), .c_out(ws0b4n1_39), .a(wand11_12), .b(wand10_13), .c_in(wand9_14));
adder_full fa142(.sum(ws0b4n0_41), .c_out(ws0b4n1_40), .a(wand10_12), .b(wand9_13), .c_in(wand8_14));
adder_full fa143(.sum(ws0b4n0_42), .c_out(ws0b4n1_41), .a(wand9_12), .b(wand8_13), .c_in(wand7_14));
adder_full fa144(.sum(ws0b4n0_43), .c_out(ws0b4n1_42), .a(wand8_12), .b(wand7_13), .c_in(wand6_14));
adder_full fa145(.sum(ws0b4n0_44), .c_out(ws0b4n1_43), .a(wand7_12), .b(wand6_13), .c_in(wand5_14));
adder_full fa146(.sum(ws0b4n0_45), .c_out(ws0b4n1_44), .a(wand6_12), .b(wand5_13), .c_in(wand4_14));
adder_full fa147(.sum(ws0b4n0_46), .c_out(ws0b4n1_45), .a(wand5_12), .b(wand4_13), .c_in(wand3_14));
adder_full fa148(.sum(ws0b4n0_47), .c_out(ws0b4n1_46), .a(wand4_12), .b(wand3_13), .c_in(wand2_14));
adder_full fa149(.sum(ws0b4n0_48), .c_out(ws0b4n1_47), .a(wand3_12), .b(wand2_13), .c_in(wand1_14));
adder_full fa150(.sum(ws0b4n0_49), .c_out(ws0b4n1_48), .a(wand2_12), .b(wand1_13), .c_in(wand0_14));
adder_half ha8(.sum(ws0b4n0_50), .c_out(ws0b4n1_49), .a(wand1_12), .b(wand0_13));
assign ws0b4n0_51 = wand0_12;
assign ws0b5n0_15 = wand31_17;
adder_half ha9(.sum(ws0b5n0_16), .c_out(ws0b5n1_15), .a(wand31_16), .b(wand30_17));
adder_full fa151(.sum(ws0b5n0_17), .c_out(ws0b5n1_16), .a(wand31_15), .b(wand30_16), .c_in(wand29_17));
adder_full fa152(.sum(ws0b5n0_18), .c_out(ws0b5n1_17), .a(wand30_15), .b(wand29_16), .c_in(wand28_17));
adder_full fa153(.sum(ws0b5n0_19), .c_out(ws0b5n1_18), .a(wand29_15), .b(wand28_16), .c_in(wand27_17));
adder_full fa154(.sum(ws0b5n0_20), .c_out(ws0b5n1_19), .a(wand28_15), .b(wand27_16), .c_in(wand26_17));
adder_full fa155(.sum(ws0b5n0_21), .c_out(ws0b5n1_20), .a(wand27_15), .b(wand26_16), .c_in(wand25_17));
adder_full fa156(.sum(ws0b5n0_22), .c_out(ws0b5n1_21), .a(wand26_15), .b(wand25_16), .c_in(wand24_17));
adder_full fa157(.sum(ws0b5n0_23), .c_out(ws0b5n1_22), .a(wand25_15), .b(wand24_16), .c_in(wand23_17));
adder_full fa158(.sum(ws0b5n0_24), .c_out(ws0b5n1_23), .a(wand24_15), .b(wand23_16), .c_in(wand22_17));
adder_full fa159(.sum(ws0b5n0_25), .c_out(ws0b5n1_24), .a(wand23_15), .b(wand22_16), .c_in(wand21_17));
adder_full fa160(.sum(ws0b5n0_26), .c_out(ws0b5n1_25), .a(wand22_15), .b(wand21_16), .c_in(wand20_17));
adder_full fa161(.sum(ws0b5n0_27), .c_out(ws0b5n1_26), .a(wand21_15), .b(wand20_16), .c_in(wand19_17));
adder_full fa162(.sum(ws0b5n0_28), .c_out(ws0b5n1_27), .a(wand20_15), .b(wand19_16), .c_in(wand18_17));
adder_full fa163(.sum(ws0b5n0_29), .c_out(ws0b5n1_28), .a(wand19_15), .b(wand18_16), .c_in(wand17_17));
adder_full fa164(.sum(ws0b5n0_30), .c_out(ws0b5n1_29), .a(wand18_15), .b(wand17_16), .c_in(wand16_17));
adder_full fa165(.sum(ws0b5n0_31), .c_out(ws0b5n1_30), .a(wand17_15), .b(wand16_16), .c_in(wand15_17));
adder_full fa166(.sum(ws0b5n0_32), .c_out(ws0b5n1_31), .a(wand16_15), .b(wand15_16), .c_in(wand14_17));
adder_full fa167(.sum(ws0b5n0_33), .c_out(ws0b5n1_32), .a(wand15_15), .b(wand14_16), .c_in(wand13_17));
adder_full fa168(.sum(ws0b5n0_34), .c_out(ws0b5n1_33), .a(wand14_15), .b(wand13_16), .c_in(wand12_17));
adder_full fa169(.sum(ws0b5n0_35), .c_out(ws0b5n1_34), .a(wand13_15), .b(wand12_16), .c_in(wand11_17));
adder_full fa170(.sum(ws0b5n0_36), .c_out(ws0b5n1_35), .a(wand12_15), .b(wand11_16), .c_in(wand10_17));
adder_full fa171(.sum(ws0b5n0_37), .c_out(ws0b5n1_36), .a(wand11_15), .b(wand10_16), .c_in(wand9_17));
adder_full fa172(.sum(ws0b5n0_38), .c_out(ws0b5n1_37), .a(wand10_15), .b(wand9_16), .c_in(wand8_17));
adder_full fa173(.sum(ws0b5n0_39), .c_out(ws0b5n1_38), .a(wand9_15), .b(wand8_16), .c_in(wand7_17));
adder_full fa174(.sum(ws0b5n0_40), .c_out(ws0b5n1_39), .a(wand8_15), .b(wand7_16), .c_in(wand6_17));
adder_full fa175(.sum(ws0b5n0_41), .c_out(ws0b5n1_40), .a(wand7_15), .b(wand6_16), .c_in(wand5_17));
adder_full fa176(.sum(ws0b5n0_42), .c_out(ws0b5n1_41), .a(wand6_15), .b(wand5_16), .c_in(wand4_17));
adder_full fa177(.sum(ws0b5n0_43), .c_out(ws0b5n1_42), .a(wand5_15), .b(wand4_16), .c_in(wand3_17));
adder_full fa178(.sum(ws0b5n0_44), .c_out(ws0b5n1_43), .a(wand4_15), .b(wand3_16), .c_in(wand2_17));
adder_full fa179(.sum(ws0b5n0_45), .c_out(ws0b5n1_44), .a(wand3_15), .b(wand2_16), .c_in(wand1_17));
adder_full fa180(.sum(ws0b5n0_46), .c_out(ws0b5n1_45), .a(wand2_15), .b(wand1_16), .c_in(wand0_17));
adder_half ha10(.sum(ws0b5n0_47), .c_out(ws0b5n1_46), .a(wand1_15), .b(wand0_16));
assign ws0b5n0_48 = wand0_15;
assign ws0b6n0_12 = wand31_20;
adder_half ha11(.sum(ws0b6n0_13), .c_out(ws0b6n1_12), .a(wand31_19), .b(wand30_20));
adder_full fa181(.sum(ws0b6n0_14), .c_out(ws0b6n1_13), .a(wand31_18), .b(wand30_19), .c_in(wand29_20));
adder_full fa182(.sum(ws0b6n0_15), .c_out(ws0b6n1_14), .a(wand30_18), .b(wand29_19), .c_in(wand28_20));
adder_full fa183(.sum(ws0b6n0_16), .c_out(ws0b6n1_15), .a(wand29_18), .b(wand28_19), .c_in(wand27_20));
adder_full fa184(.sum(ws0b6n0_17), .c_out(ws0b6n1_16), .a(wand28_18), .b(wand27_19), .c_in(wand26_20));
adder_full fa185(.sum(ws0b6n0_18), .c_out(ws0b6n1_17), .a(wand27_18), .b(wand26_19), .c_in(wand25_20));
adder_full fa186(.sum(ws0b6n0_19), .c_out(ws0b6n1_18), .a(wand26_18), .b(wand25_19), .c_in(wand24_20));
adder_full fa187(.sum(ws0b6n0_20), .c_out(ws0b6n1_19), .a(wand25_18), .b(wand24_19), .c_in(wand23_20));
adder_full fa188(.sum(ws0b6n0_21), .c_out(ws0b6n1_20), .a(wand24_18), .b(wand23_19), .c_in(wand22_20));
adder_full fa189(.sum(ws0b6n0_22), .c_out(ws0b6n1_21), .a(wand23_18), .b(wand22_19), .c_in(wand21_20));
adder_full fa190(.sum(ws0b6n0_23), .c_out(ws0b6n1_22), .a(wand22_18), .b(wand21_19), .c_in(wand20_20));
adder_full fa191(.sum(ws0b6n0_24), .c_out(ws0b6n1_23), .a(wand21_18), .b(wand20_19), .c_in(wand19_20));
adder_full fa192(.sum(ws0b6n0_25), .c_out(ws0b6n1_24), .a(wand20_18), .b(wand19_19), .c_in(wand18_20));
adder_full fa193(.sum(ws0b6n0_26), .c_out(ws0b6n1_25), .a(wand19_18), .b(wand18_19), .c_in(wand17_20));
adder_full fa194(.sum(ws0b6n0_27), .c_out(ws0b6n1_26), .a(wand18_18), .b(wand17_19), .c_in(wand16_20));
adder_full fa195(.sum(ws0b6n0_28), .c_out(ws0b6n1_27), .a(wand17_18), .b(wand16_19), .c_in(wand15_20));
adder_full fa196(.sum(ws0b6n0_29), .c_out(ws0b6n1_28), .a(wand16_18), .b(wand15_19), .c_in(wand14_20));
adder_full fa197(.sum(ws0b6n0_30), .c_out(ws0b6n1_29), .a(wand15_18), .b(wand14_19), .c_in(wand13_20));
adder_full fa198(.sum(ws0b6n0_31), .c_out(ws0b6n1_30), .a(wand14_18), .b(wand13_19), .c_in(wand12_20));
adder_full fa199(.sum(ws0b6n0_32), .c_out(ws0b6n1_31), .a(wand13_18), .b(wand12_19), .c_in(wand11_20));
adder_full fa200(.sum(ws0b6n0_33), .c_out(ws0b6n1_32), .a(wand12_18), .b(wand11_19), .c_in(wand10_20));
adder_full fa201(.sum(ws0b6n0_34), .c_out(ws0b6n1_33), .a(wand11_18), .b(wand10_19), .c_in(wand9_20));
adder_full fa202(.sum(ws0b6n0_35), .c_out(ws0b6n1_34), .a(wand10_18), .b(wand9_19), .c_in(wand8_20));
adder_full fa203(.sum(ws0b6n0_36), .c_out(ws0b6n1_35), .a(wand9_18), .b(wand8_19), .c_in(wand7_20));
adder_full fa204(.sum(ws0b6n0_37), .c_out(ws0b6n1_36), .a(wand8_18), .b(wand7_19), .c_in(wand6_20));
adder_full fa205(.sum(ws0b6n0_38), .c_out(ws0b6n1_37), .a(wand7_18), .b(wand6_19), .c_in(wand5_20));
adder_full fa206(.sum(ws0b6n0_39), .c_out(ws0b6n1_38), .a(wand6_18), .b(wand5_19), .c_in(wand4_20));
adder_full fa207(.sum(ws0b6n0_40), .c_out(ws0b6n1_39), .a(wand5_18), .b(wand4_19), .c_in(wand3_20));
adder_full fa208(.sum(ws0b6n0_41), .c_out(ws0b6n1_40), .a(wand4_18), .b(wand3_19), .c_in(wand2_20));
adder_full fa209(.sum(ws0b6n0_42), .c_out(ws0b6n1_41), .a(wand3_18), .b(wand2_19), .c_in(wand1_20));
adder_full fa210(.sum(ws0b6n0_43), .c_out(ws0b6n1_42), .a(wand2_18), .b(wand1_19), .c_in(wand0_20));
adder_half ha12(.sum(ws0b6n0_44), .c_out(ws0b6n1_43), .a(wand1_18), .b(wand0_19));
assign ws0b6n0_45 = wand0_18;
assign ws0b7n0_9 = wand31_23;
adder_half ha13(.sum(ws0b7n0_10), .c_out(ws0b7n1_9), .a(wand31_22), .b(wand30_23));
adder_full fa211(.sum(ws0b7n0_11), .c_out(ws0b7n1_10), .a(wand31_21), .b(wand30_22), .c_in(wand29_23));
adder_full fa212(.sum(ws0b7n0_12), .c_out(ws0b7n1_11), .a(wand30_21), .b(wand29_22), .c_in(wand28_23));
adder_full fa213(.sum(ws0b7n0_13), .c_out(ws0b7n1_12), .a(wand29_21), .b(wand28_22), .c_in(wand27_23));
adder_full fa214(.sum(ws0b7n0_14), .c_out(ws0b7n1_13), .a(wand28_21), .b(wand27_22), .c_in(wand26_23));
adder_full fa215(.sum(ws0b7n0_15), .c_out(ws0b7n1_14), .a(wand27_21), .b(wand26_22), .c_in(wand25_23));
adder_full fa216(.sum(ws0b7n0_16), .c_out(ws0b7n1_15), .a(wand26_21), .b(wand25_22), .c_in(wand24_23));
adder_full fa217(.sum(ws0b7n0_17), .c_out(ws0b7n1_16), .a(wand25_21), .b(wand24_22), .c_in(wand23_23));
adder_full fa218(.sum(ws0b7n0_18), .c_out(ws0b7n1_17), .a(wand24_21), .b(wand23_22), .c_in(wand22_23));
adder_full fa219(.sum(ws0b7n0_19), .c_out(ws0b7n1_18), .a(wand23_21), .b(wand22_22), .c_in(wand21_23));
adder_full fa220(.sum(ws0b7n0_20), .c_out(ws0b7n1_19), .a(wand22_21), .b(wand21_22), .c_in(wand20_23));
adder_full fa221(.sum(ws0b7n0_21), .c_out(ws0b7n1_20), .a(wand21_21), .b(wand20_22), .c_in(wand19_23));
adder_full fa222(.sum(ws0b7n0_22), .c_out(ws0b7n1_21), .a(wand20_21), .b(wand19_22), .c_in(wand18_23));
adder_full fa223(.sum(ws0b7n0_23), .c_out(ws0b7n1_22), .a(wand19_21), .b(wand18_22), .c_in(wand17_23));
adder_full fa224(.sum(ws0b7n0_24), .c_out(ws0b7n1_23), .a(wand18_21), .b(wand17_22), .c_in(wand16_23));
adder_full fa225(.sum(ws0b7n0_25), .c_out(ws0b7n1_24), .a(wand17_21), .b(wand16_22), .c_in(wand15_23));
adder_full fa226(.sum(ws0b7n0_26), .c_out(ws0b7n1_25), .a(wand16_21), .b(wand15_22), .c_in(wand14_23));
adder_full fa227(.sum(ws0b7n0_27), .c_out(ws0b7n1_26), .a(wand15_21), .b(wand14_22), .c_in(wand13_23));
adder_full fa228(.sum(ws0b7n0_28), .c_out(ws0b7n1_27), .a(wand14_21), .b(wand13_22), .c_in(wand12_23));
adder_full fa229(.sum(ws0b7n0_29), .c_out(ws0b7n1_28), .a(wand13_21), .b(wand12_22), .c_in(wand11_23));
adder_full fa230(.sum(ws0b7n0_30), .c_out(ws0b7n1_29), .a(wand12_21), .b(wand11_22), .c_in(wand10_23));
adder_full fa231(.sum(ws0b7n0_31), .c_out(ws0b7n1_30), .a(wand11_21), .b(wand10_22), .c_in(wand9_23));
adder_full fa232(.sum(ws0b7n0_32), .c_out(ws0b7n1_31), .a(wand10_21), .b(wand9_22), .c_in(wand8_23));
adder_full fa233(.sum(ws0b7n0_33), .c_out(ws0b7n1_32), .a(wand9_21), .b(wand8_22), .c_in(wand7_23));
adder_full fa234(.sum(ws0b7n0_34), .c_out(ws0b7n1_33), .a(wand8_21), .b(wand7_22), .c_in(wand6_23));
adder_full fa235(.sum(ws0b7n0_35), .c_out(ws0b7n1_34), .a(wand7_21), .b(wand6_22), .c_in(wand5_23));
adder_full fa236(.sum(ws0b7n0_36), .c_out(ws0b7n1_35), .a(wand6_21), .b(wand5_22), .c_in(wand4_23));
adder_full fa237(.sum(ws0b7n0_37), .c_out(ws0b7n1_36), .a(wand5_21), .b(wand4_22), .c_in(wand3_23));
adder_full fa238(.sum(ws0b7n0_38), .c_out(ws0b7n1_37), .a(wand4_21), .b(wand3_22), .c_in(wand2_23));
adder_full fa239(.sum(ws0b7n0_39), .c_out(ws0b7n1_38), .a(wand3_21), .b(wand2_22), .c_in(wand1_23));
adder_full fa240(.sum(ws0b7n0_40), .c_out(ws0b7n1_39), .a(wand2_21), .b(wand1_22), .c_in(wand0_23));
adder_half ha14(.sum(ws0b7n0_41), .c_out(ws0b7n1_40), .a(wand1_21), .b(wand0_22));
assign ws0b7n0_42 = wand0_21;
assign ws0b8n0_6 = wand31_26;
adder_half ha15(.sum(ws0b8n0_7), .c_out(ws0b8n1_6), .a(wand31_25), .b(wand30_26));
adder_full fa241(.sum(ws0b8n0_8), .c_out(ws0b8n1_7), .a(wand31_24), .b(wand30_25), .c_in(wand29_26));
adder_full fa242(.sum(ws0b8n0_9), .c_out(ws0b8n1_8), .a(wand30_24), .b(wand29_25), .c_in(wand28_26));
adder_full fa243(.sum(ws0b8n0_10), .c_out(ws0b8n1_9), .a(wand29_24), .b(wand28_25), .c_in(wand27_26));
adder_full fa244(.sum(ws0b8n0_11), .c_out(ws0b8n1_10), .a(wand28_24), .b(wand27_25), .c_in(wand26_26));
adder_full fa245(.sum(ws0b8n0_12), .c_out(ws0b8n1_11), .a(wand27_24), .b(wand26_25), .c_in(wand25_26));
adder_full fa246(.sum(ws0b8n0_13), .c_out(ws0b8n1_12), .a(wand26_24), .b(wand25_25), .c_in(wand24_26));
adder_full fa247(.sum(ws0b8n0_14), .c_out(ws0b8n1_13), .a(wand25_24), .b(wand24_25), .c_in(wand23_26));
adder_full fa248(.sum(ws0b8n0_15), .c_out(ws0b8n1_14), .a(wand24_24), .b(wand23_25), .c_in(wand22_26));
adder_full fa249(.sum(ws0b8n0_16), .c_out(ws0b8n1_15), .a(wand23_24), .b(wand22_25), .c_in(wand21_26));
adder_full fa250(.sum(ws0b8n0_17), .c_out(ws0b8n1_16), .a(wand22_24), .b(wand21_25), .c_in(wand20_26));
adder_full fa251(.sum(ws0b8n0_18), .c_out(ws0b8n1_17), .a(wand21_24), .b(wand20_25), .c_in(wand19_26));
adder_full fa252(.sum(ws0b8n0_19), .c_out(ws0b8n1_18), .a(wand20_24), .b(wand19_25), .c_in(wand18_26));
adder_full fa253(.sum(ws0b8n0_20), .c_out(ws0b8n1_19), .a(wand19_24), .b(wand18_25), .c_in(wand17_26));
adder_full fa254(.sum(ws0b8n0_21), .c_out(ws0b8n1_20), .a(wand18_24), .b(wand17_25), .c_in(wand16_26));
adder_full fa255(.sum(ws0b8n0_22), .c_out(ws0b8n1_21), .a(wand17_24), .b(wand16_25), .c_in(wand15_26));
adder_full fa256(.sum(ws0b8n0_23), .c_out(ws0b8n1_22), .a(wand16_24), .b(wand15_25), .c_in(wand14_26));
adder_full fa257(.sum(ws0b8n0_24), .c_out(ws0b8n1_23), .a(wand15_24), .b(wand14_25), .c_in(wand13_26));
adder_full fa258(.sum(ws0b8n0_25), .c_out(ws0b8n1_24), .a(wand14_24), .b(wand13_25), .c_in(wand12_26));
adder_full fa259(.sum(ws0b8n0_26), .c_out(ws0b8n1_25), .a(wand13_24), .b(wand12_25), .c_in(wand11_26));
adder_full fa260(.sum(ws0b8n0_27), .c_out(ws0b8n1_26), .a(wand12_24), .b(wand11_25), .c_in(wand10_26));
adder_full fa261(.sum(ws0b8n0_28), .c_out(ws0b8n1_27), .a(wand11_24), .b(wand10_25), .c_in(wand9_26));
adder_full fa262(.sum(ws0b8n0_29), .c_out(ws0b8n1_28), .a(wand10_24), .b(wand9_25), .c_in(wand8_26));
adder_full fa263(.sum(ws0b8n0_30), .c_out(ws0b8n1_29), .a(wand9_24), .b(wand8_25), .c_in(wand7_26));
adder_full fa264(.sum(ws0b8n0_31), .c_out(ws0b8n1_30), .a(wand8_24), .b(wand7_25), .c_in(wand6_26));
adder_full fa265(.sum(ws0b8n0_32), .c_out(ws0b8n1_31), .a(wand7_24), .b(wand6_25), .c_in(wand5_26));
adder_full fa266(.sum(ws0b8n0_33), .c_out(ws0b8n1_32), .a(wand6_24), .b(wand5_25), .c_in(wand4_26));
adder_full fa267(.sum(ws0b8n0_34), .c_out(ws0b8n1_33), .a(wand5_24), .b(wand4_25), .c_in(wand3_26));
adder_full fa268(.sum(ws0b8n0_35), .c_out(ws0b8n1_34), .a(wand4_24), .b(wand3_25), .c_in(wand2_26));
adder_full fa269(.sum(ws0b8n0_36), .c_out(ws0b8n1_35), .a(wand3_24), .b(wand2_25), .c_in(wand1_26));
adder_full fa270(.sum(ws0b8n0_37), .c_out(ws0b8n1_36), .a(wand2_24), .b(wand1_25), .c_in(wand0_26));
adder_half ha16(.sum(ws0b8n0_38), .c_out(ws0b8n1_37), .a(wand1_24), .b(wand0_25));
assign ws0b8n0_39 = wand0_24;
assign ws0b9n0_3 = wand31_29;
adder_half ha17(.sum(ws0b9n0_4), .c_out(ws0b9n1_3), .a(wand31_28), .b(wand30_29));
adder_full fa271(.sum(ws0b9n0_5), .c_out(ws0b9n1_4), .a(wand31_27), .b(wand30_28), .c_in(wand29_29));
adder_full fa272(.sum(ws0b9n0_6), .c_out(ws0b9n1_5), .a(wand30_27), .b(wand29_28), .c_in(wand28_29));
adder_full fa273(.sum(ws0b9n0_7), .c_out(ws0b9n1_6), .a(wand29_27), .b(wand28_28), .c_in(wand27_29));
adder_full fa274(.sum(ws0b9n0_8), .c_out(ws0b9n1_7), .a(wand28_27), .b(wand27_28), .c_in(wand26_29));
adder_full fa275(.sum(ws0b9n0_9), .c_out(ws0b9n1_8), .a(wand27_27), .b(wand26_28), .c_in(wand25_29));
adder_full fa276(.sum(ws0b9n0_10), .c_out(ws0b9n1_9), .a(wand26_27), .b(wand25_28), .c_in(wand24_29));
adder_full fa277(.sum(ws0b9n0_11), .c_out(ws0b9n1_10), .a(wand25_27), .b(wand24_28), .c_in(wand23_29));
adder_full fa278(.sum(ws0b9n0_12), .c_out(ws0b9n1_11), .a(wand24_27), .b(wand23_28), .c_in(wand22_29));
adder_full fa279(.sum(ws0b9n0_13), .c_out(ws0b9n1_12), .a(wand23_27), .b(wand22_28), .c_in(wand21_29));
adder_full fa280(.sum(ws0b9n0_14), .c_out(ws0b9n1_13), .a(wand22_27), .b(wand21_28), .c_in(wand20_29));
adder_full fa281(.sum(ws0b9n0_15), .c_out(ws0b9n1_14), .a(wand21_27), .b(wand20_28), .c_in(wand19_29));
adder_full fa282(.sum(ws0b9n0_16), .c_out(ws0b9n1_15), .a(wand20_27), .b(wand19_28), .c_in(wand18_29));
adder_full fa283(.sum(ws0b9n0_17), .c_out(ws0b9n1_16), .a(wand19_27), .b(wand18_28), .c_in(wand17_29));
adder_full fa284(.sum(ws0b9n0_18), .c_out(ws0b9n1_17), .a(wand18_27), .b(wand17_28), .c_in(wand16_29));
adder_full fa285(.sum(ws0b9n0_19), .c_out(ws0b9n1_18), .a(wand17_27), .b(wand16_28), .c_in(wand15_29));
adder_full fa286(.sum(ws0b9n0_20), .c_out(ws0b9n1_19), .a(wand16_27), .b(wand15_28), .c_in(wand14_29));
adder_full fa287(.sum(ws0b9n0_21), .c_out(ws0b9n1_20), .a(wand15_27), .b(wand14_28), .c_in(wand13_29));
adder_full fa288(.sum(ws0b9n0_22), .c_out(ws0b9n1_21), .a(wand14_27), .b(wand13_28), .c_in(wand12_29));
adder_full fa289(.sum(ws0b9n0_23), .c_out(ws0b9n1_22), .a(wand13_27), .b(wand12_28), .c_in(wand11_29));
adder_full fa290(.sum(ws0b9n0_24), .c_out(ws0b9n1_23), .a(wand12_27), .b(wand11_28), .c_in(wand10_29));
adder_full fa291(.sum(ws0b9n0_25), .c_out(ws0b9n1_24), .a(wand11_27), .b(wand10_28), .c_in(wand9_29));
adder_full fa292(.sum(ws0b9n0_26), .c_out(ws0b9n1_25), .a(wand10_27), .b(wand9_28), .c_in(wand8_29));
adder_full fa293(.sum(ws0b9n0_27), .c_out(ws0b9n1_26), .a(wand9_27), .b(wand8_28), .c_in(wand7_29));
adder_full fa294(.sum(ws0b9n0_28), .c_out(ws0b9n1_27), .a(wand8_27), .b(wand7_28), .c_in(wand6_29));
adder_full fa295(.sum(ws0b9n0_29), .c_out(ws0b9n1_28), .a(wand7_27), .b(wand6_28), .c_in(wand5_29));
adder_full fa296(.sum(ws0b9n0_30), .c_out(ws0b9n1_29), .a(wand6_27), .b(wand5_28), .c_in(wand4_29));
adder_full fa297(.sum(ws0b9n0_31), .c_out(ws0b9n1_30), .a(wand5_27), .b(wand4_28), .c_in(wand3_29));
adder_full fa298(.sum(ws0b9n0_32), .c_out(ws0b9n1_31), .a(wand4_27), .b(wand3_28), .c_in(wand2_29));
adder_full fa299(.sum(ws0b9n0_33), .c_out(ws0b9n1_32), .a(wand3_27), .b(wand2_28), .c_in(wand1_29));
adder_full fa300(.sum(ws0b9n0_34), .c_out(ws0b9n1_33), .a(wand2_27), .b(wand1_28), .c_in(wand0_29));
adder_half ha18(.sum(ws0b9n0_35), .c_out(ws0b9n1_34), .a(wand1_27), .b(wand0_28));
assign ws0b9n0_36 = wand0_27;

assign ws1b0n0_27 = ws0b1n0_27;
assign ws1b0n0_28 = ws0b1n0_28;
assign ws1b0n0_29 = ws0b1n0_29;
adder_full fa301(.sum(ws1b0n0_30), .c_out(ws1b0n1_29), .a(ws0b0n0_30), .b(ws0b0n1_30), .c_in(ws0b1n0_30));
adder_full fa302(.sum(ws1b0n0_31), .c_out(ws1b0n1_30), .a(ws0b0n0_31), .b(ws0b0n1_31), .c_in(ws0b1n0_31));
adder_full fa303(.sum(ws1b0n0_32), .c_out(ws1b0n1_31), .a(ws0b0n0_32), .b(ws0b0n1_32), .c_in(ws0b1n0_32));
adder_full fa304(.sum(ws1b0n0_33), .c_out(ws1b0n1_32), .a(ws0b0n0_33), .b(ws0b0n1_33), .c_in(ws0b1n0_33));
adder_full fa305(.sum(ws1b0n0_34), .c_out(ws1b0n1_33), .a(ws0b0n0_34), .b(ws0b0n1_34), .c_in(ws0b1n0_34));
adder_full fa306(.sum(ws1b0n0_35), .c_out(ws1b0n1_34), .a(ws0b0n0_35), .b(ws0b0n1_35), .c_in(ws0b1n0_35));
adder_full fa307(.sum(ws1b0n0_36), .c_out(ws1b0n1_35), .a(ws0b0n0_36), .b(ws0b0n1_36), .c_in(ws0b1n0_36));
adder_full fa308(.sum(ws1b0n0_37), .c_out(ws1b0n1_36), .a(ws0b0n0_37), .b(ws0b0n1_37), .c_in(ws0b1n0_37));
adder_full fa309(.sum(ws1b0n0_38), .c_out(ws1b0n1_37), .a(ws0b0n0_38), .b(ws0b0n1_38), .c_in(ws0b1n0_38));
adder_full fa310(.sum(ws1b0n0_39), .c_out(ws1b0n1_38), .a(ws0b0n0_39), .b(ws0b0n1_39), .c_in(ws0b1n0_39));
adder_full fa311(.sum(ws1b0n0_40), .c_out(ws1b0n1_39), .a(ws0b0n0_40), .b(ws0b0n1_40), .c_in(ws0b1n0_40));
adder_full fa312(.sum(ws1b0n0_41), .c_out(ws1b0n1_40), .a(ws0b0n0_41), .b(ws0b0n1_41), .c_in(ws0b1n0_41));
adder_full fa313(.sum(ws1b0n0_42), .c_out(ws1b0n1_41), .a(ws0b0n0_42), .b(ws0b0n1_42), .c_in(ws0b1n0_42));
adder_full fa314(.sum(ws1b0n0_43), .c_out(ws1b0n1_42), .a(ws0b0n0_43), .b(ws0b0n1_43), .c_in(ws0b1n0_43));
adder_full fa315(.sum(ws1b0n0_44), .c_out(ws1b0n1_43), .a(ws0b0n0_44), .b(ws0b0n1_44), .c_in(ws0b1n0_44));
adder_full fa316(.sum(ws1b0n0_45), .c_out(ws1b0n1_44), .a(ws0b0n0_45), .b(ws0b0n1_45), .c_in(ws0b1n0_45));
adder_full fa317(.sum(ws1b0n0_46), .c_out(ws1b0n1_45), .a(ws0b0n0_46), .b(ws0b0n1_46), .c_in(ws0b1n0_46));
adder_full fa318(.sum(ws1b0n0_47), .c_out(ws1b0n1_46), .a(ws0b0n0_47), .b(ws0b0n1_47), .c_in(ws0b1n0_47));
adder_full fa319(.sum(ws1b0n0_48), .c_out(ws1b0n1_47), .a(ws0b0n0_48), .b(ws0b0n1_48), .c_in(ws0b1n0_48));
adder_full fa320(.sum(ws1b0n0_49), .c_out(ws1b0n1_48), .a(ws0b0n0_49), .b(ws0b0n1_49), .c_in(ws0b1n0_49));
adder_full fa321(.sum(ws1b0n0_50), .c_out(ws1b0n1_49), .a(ws0b0n0_50), .b(ws0b0n1_50), .c_in(ws0b1n0_50));
adder_full fa322(.sum(ws1b0n0_51), .c_out(ws1b0n1_50), .a(ws0b0n0_51), .b(ws0b0n1_51), .c_in(ws0b1n0_51));
adder_full fa323(.sum(ws1b0n0_52), .c_out(ws1b0n1_51), .a(ws0b0n0_52), .b(ws0b0n1_52), .c_in(ws0b1n0_52));
adder_full fa324(.sum(ws1b0n0_53), .c_out(ws1b0n1_52), .a(ws0b0n0_53), .b(ws0b0n1_53), .c_in(ws0b1n0_53));
adder_full fa325(.sum(ws1b0n0_54), .c_out(ws1b0n1_53), .a(ws0b0n0_54), .b(ws0b0n1_54), .c_in(ws0b1n0_54));
adder_full fa326(.sum(ws1b0n0_55), .c_out(ws1b0n1_54), .a(ws0b0n0_55), .b(ws0b0n1_55), .c_in(ws0b1n0_55));
adder_full fa327(.sum(ws1b0n0_56), .c_out(ws1b0n1_55), .a(ws0b0n0_56), .b(ws0b0n1_56), .c_in(ws0b1n0_56));
adder_full fa328(.sum(ws1b0n0_57), .c_out(ws1b0n1_56), .a(ws0b0n0_57), .b(ws0b0n1_57), .c_in(ws0b1n0_57));
adder_full fa329(.sum(ws1b0n0_58), .c_out(ws1b0n1_57), .a(ws0b0n0_58), .b(ws0b0n1_58), .c_in(ws0b1n0_58));
adder_full fa330(.sum(ws1b0n0_59), .c_out(ws1b0n1_58), .a(ws0b0n0_59), .b(ws0b0n1_59), .c_in(ws0b1n0_59));
adder_full fa331(.sum(ws1b0n0_60), .c_out(ws1b0n1_59), .a(ws0b0n0_60), .b(ws0b0n1_60), .c_in(ws0b1n0_60));
adder_half ha19(.sum(ws1b0n0_61), .c_out(ws1b0n1_60), .a(ws0b0n0_61), .b(ws0b0n1_61));
assign ws1b0n0_62 = ws0b0n0_62;
assign ws1b0n0_63 = ws0b0n0_63;
adder_half ha20(.sum(ws1b1n0_24), .c_out(ws1b1n1_23), .a(ws0b2n0_24), .b(ws0b2n1_24));
adder_half ha21(.sum(ws1b1n0_25), .c_out(ws1b1n1_24), .a(ws0b2n0_25), .b(ws0b2n1_25));
adder_half ha22(.sum(ws1b1n0_26), .c_out(ws1b1n1_25), .a(ws0b2n0_26), .b(ws0b2n1_26));
adder_full fa332(.sum(ws1b1n0_27), .c_out(ws1b1n1_26), .a(ws0b1n1_27), .b(ws0b2n0_27), .c_in(ws0b2n1_27));
adder_full fa333(.sum(ws1b1n0_28), .c_out(ws1b1n1_27), .a(ws0b1n1_28), .b(ws0b2n0_28), .c_in(ws0b2n1_28));
adder_full fa334(.sum(ws1b1n0_29), .c_out(ws1b1n1_28), .a(ws0b1n1_29), .b(ws0b2n0_29), .c_in(ws0b2n1_29));
adder_full fa335(.sum(ws1b1n0_30), .c_out(ws1b1n1_29), .a(ws0b1n1_30), .b(ws0b2n0_30), .c_in(ws0b2n1_30));
adder_full fa336(.sum(ws1b1n0_31), .c_out(ws1b1n1_30), .a(ws0b1n1_31), .b(ws0b2n0_31), .c_in(ws0b2n1_31));
adder_full fa337(.sum(ws1b1n0_32), .c_out(ws1b1n1_31), .a(ws0b1n1_32), .b(ws0b2n0_32), .c_in(ws0b2n1_32));
adder_full fa338(.sum(ws1b1n0_33), .c_out(ws1b1n1_32), .a(ws0b1n1_33), .b(ws0b2n0_33), .c_in(ws0b2n1_33));
adder_full fa339(.sum(ws1b1n0_34), .c_out(ws1b1n1_33), .a(ws0b1n1_34), .b(ws0b2n0_34), .c_in(ws0b2n1_34));
adder_full fa340(.sum(ws1b1n0_35), .c_out(ws1b1n1_34), .a(ws0b1n1_35), .b(ws0b2n0_35), .c_in(ws0b2n1_35));
adder_full fa341(.sum(ws1b1n0_36), .c_out(ws1b1n1_35), .a(ws0b1n1_36), .b(ws0b2n0_36), .c_in(ws0b2n1_36));
adder_full fa342(.sum(ws1b1n0_37), .c_out(ws1b1n1_36), .a(ws0b1n1_37), .b(ws0b2n0_37), .c_in(ws0b2n1_37));
adder_full fa343(.sum(ws1b1n0_38), .c_out(ws1b1n1_37), .a(ws0b1n1_38), .b(ws0b2n0_38), .c_in(ws0b2n1_38));
adder_full fa344(.sum(ws1b1n0_39), .c_out(ws1b1n1_38), .a(ws0b1n1_39), .b(ws0b2n0_39), .c_in(ws0b2n1_39));
adder_full fa345(.sum(ws1b1n0_40), .c_out(ws1b1n1_39), .a(ws0b1n1_40), .b(ws0b2n0_40), .c_in(ws0b2n1_40));
adder_full fa346(.sum(ws1b1n0_41), .c_out(ws1b1n1_40), .a(ws0b1n1_41), .b(ws0b2n0_41), .c_in(ws0b2n1_41));
adder_full fa347(.sum(ws1b1n0_42), .c_out(ws1b1n1_41), .a(ws0b1n1_42), .b(ws0b2n0_42), .c_in(ws0b2n1_42));
adder_full fa348(.sum(ws1b1n0_43), .c_out(ws1b1n1_42), .a(ws0b1n1_43), .b(ws0b2n0_43), .c_in(ws0b2n1_43));
adder_full fa349(.sum(ws1b1n0_44), .c_out(ws1b1n1_43), .a(ws0b1n1_44), .b(ws0b2n0_44), .c_in(ws0b2n1_44));
adder_full fa350(.sum(ws1b1n0_45), .c_out(ws1b1n1_44), .a(ws0b1n1_45), .b(ws0b2n0_45), .c_in(ws0b2n1_45));
adder_full fa351(.sum(ws1b1n0_46), .c_out(ws1b1n1_45), .a(ws0b1n1_46), .b(ws0b2n0_46), .c_in(ws0b2n1_46));
adder_full fa352(.sum(ws1b1n0_47), .c_out(ws1b1n1_46), .a(ws0b1n1_47), .b(ws0b2n0_47), .c_in(ws0b2n1_47));
adder_full fa353(.sum(ws1b1n0_48), .c_out(ws1b1n1_47), .a(ws0b1n1_48), .b(ws0b2n0_48), .c_in(ws0b2n1_48));
adder_full fa354(.sum(ws1b1n0_49), .c_out(ws1b1n1_48), .a(ws0b1n1_49), .b(ws0b2n0_49), .c_in(ws0b2n1_49));
adder_full fa355(.sum(ws1b1n0_50), .c_out(ws1b1n1_49), .a(ws0b1n1_50), .b(ws0b2n0_50), .c_in(ws0b2n1_50));
adder_full fa356(.sum(ws1b1n0_51), .c_out(ws1b1n1_50), .a(ws0b1n1_51), .b(ws0b2n0_51), .c_in(ws0b2n1_51));
adder_full fa357(.sum(ws1b1n0_52), .c_out(ws1b1n1_51), .a(ws0b1n1_52), .b(ws0b2n0_52), .c_in(ws0b2n1_52));
adder_full fa358(.sum(ws1b1n0_53), .c_out(ws1b1n1_52), .a(ws0b1n1_53), .b(ws0b2n0_53), .c_in(ws0b2n1_53));
adder_full fa359(.sum(ws1b1n0_54), .c_out(ws1b1n1_53), .a(ws0b1n1_54), .b(ws0b2n0_54), .c_in(ws0b2n1_54));
adder_full fa360(.sum(ws1b1n0_55), .c_out(ws1b1n1_54), .a(ws0b1n1_55), .b(ws0b2n0_55), .c_in(ws0b2n1_55));
adder_half ha23(.sum(ws1b1n0_56), .c_out(ws1b1n1_55), .a(ws0b1n1_56), .b(ws0b2n0_56));
adder_half ha24(.sum(ws1b1n0_57), .c_out(ws1b1n1_56), .a(ws0b1n1_57), .b(ws0b2n0_57));
assign ws1b1n0_58 = ws0b1n1_58;
assign ws1b2n0_18 = ws0b4n0_18;
assign ws1b2n0_19 = ws0b4n0_19;
assign ws1b2n0_20 = ws0b4n0_20;
adder_full fa361(.sum(ws1b2n0_21), .c_out(ws1b2n1_20), .a(ws0b3n0_21), .b(ws0b3n1_21), .c_in(ws0b4n0_21));
adder_full fa362(.sum(ws1b2n0_22), .c_out(ws1b2n1_21), .a(ws0b3n0_22), .b(ws0b3n1_22), .c_in(ws0b4n0_22));
adder_full fa363(.sum(ws1b2n0_23), .c_out(ws1b2n1_22), .a(ws0b3n0_23), .b(ws0b3n1_23), .c_in(ws0b4n0_23));
adder_full fa364(.sum(ws1b2n0_24), .c_out(ws1b2n1_23), .a(ws0b3n0_24), .b(ws0b3n1_24), .c_in(ws0b4n0_24));
adder_full fa365(.sum(ws1b2n0_25), .c_out(ws1b2n1_24), .a(ws0b3n0_25), .b(ws0b3n1_25), .c_in(ws0b4n0_25));
adder_full fa366(.sum(ws1b2n0_26), .c_out(ws1b2n1_25), .a(ws0b3n0_26), .b(ws0b3n1_26), .c_in(ws0b4n0_26));
adder_full fa367(.sum(ws1b2n0_27), .c_out(ws1b2n1_26), .a(ws0b3n0_27), .b(ws0b3n1_27), .c_in(ws0b4n0_27));
adder_full fa368(.sum(ws1b2n0_28), .c_out(ws1b2n1_27), .a(ws0b3n0_28), .b(ws0b3n1_28), .c_in(ws0b4n0_28));
adder_full fa369(.sum(ws1b2n0_29), .c_out(ws1b2n1_28), .a(ws0b3n0_29), .b(ws0b3n1_29), .c_in(ws0b4n0_29));
adder_full fa370(.sum(ws1b2n0_30), .c_out(ws1b2n1_29), .a(ws0b3n0_30), .b(ws0b3n1_30), .c_in(ws0b4n0_30));
adder_full fa371(.sum(ws1b2n0_31), .c_out(ws1b2n1_30), .a(ws0b3n0_31), .b(ws0b3n1_31), .c_in(ws0b4n0_31));
adder_full fa372(.sum(ws1b2n0_32), .c_out(ws1b2n1_31), .a(ws0b3n0_32), .b(ws0b3n1_32), .c_in(ws0b4n0_32));
adder_full fa373(.sum(ws1b2n0_33), .c_out(ws1b2n1_32), .a(ws0b3n0_33), .b(ws0b3n1_33), .c_in(ws0b4n0_33));
adder_full fa374(.sum(ws1b2n0_34), .c_out(ws1b2n1_33), .a(ws0b3n0_34), .b(ws0b3n1_34), .c_in(ws0b4n0_34));
adder_full fa375(.sum(ws1b2n0_35), .c_out(ws1b2n1_34), .a(ws0b3n0_35), .b(ws0b3n1_35), .c_in(ws0b4n0_35));
adder_full fa376(.sum(ws1b2n0_36), .c_out(ws1b2n1_35), .a(ws0b3n0_36), .b(ws0b3n1_36), .c_in(ws0b4n0_36));
adder_full fa377(.sum(ws1b2n0_37), .c_out(ws1b2n1_36), .a(ws0b3n0_37), .b(ws0b3n1_37), .c_in(ws0b4n0_37));
adder_full fa378(.sum(ws1b2n0_38), .c_out(ws1b2n1_37), .a(ws0b3n0_38), .b(ws0b3n1_38), .c_in(ws0b4n0_38));
adder_full fa379(.sum(ws1b2n0_39), .c_out(ws1b2n1_38), .a(ws0b3n0_39), .b(ws0b3n1_39), .c_in(ws0b4n0_39));
adder_full fa380(.sum(ws1b2n0_40), .c_out(ws1b2n1_39), .a(ws0b3n0_40), .b(ws0b3n1_40), .c_in(ws0b4n0_40));
adder_full fa381(.sum(ws1b2n0_41), .c_out(ws1b2n1_40), .a(ws0b3n0_41), .b(ws0b3n1_41), .c_in(ws0b4n0_41));
adder_full fa382(.sum(ws1b2n0_42), .c_out(ws1b2n1_41), .a(ws0b3n0_42), .b(ws0b3n1_42), .c_in(ws0b4n0_42));
adder_full fa383(.sum(ws1b2n0_43), .c_out(ws1b2n1_42), .a(ws0b3n0_43), .b(ws0b3n1_43), .c_in(ws0b4n0_43));
adder_full fa384(.sum(ws1b2n0_44), .c_out(ws1b2n1_43), .a(ws0b3n0_44), .b(ws0b3n1_44), .c_in(ws0b4n0_44));
adder_full fa385(.sum(ws1b2n0_45), .c_out(ws1b2n1_44), .a(ws0b3n0_45), .b(ws0b3n1_45), .c_in(ws0b4n0_45));
adder_full fa386(.sum(ws1b2n0_46), .c_out(ws1b2n1_45), .a(ws0b3n0_46), .b(ws0b3n1_46), .c_in(ws0b4n0_46));
adder_full fa387(.sum(ws1b2n0_47), .c_out(ws1b2n1_46), .a(ws0b3n0_47), .b(ws0b3n1_47), .c_in(ws0b4n0_47));
adder_full fa388(.sum(ws1b2n0_48), .c_out(ws1b2n1_47), .a(ws0b3n0_48), .b(ws0b3n1_48), .c_in(ws0b4n0_48));
adder_full fa389(.sum(ws1b2n0_49), .c_out(ws1b2n1_48), .a(ws0b3n0_49), .b(ws0b3n1_49), .c_in(ws0b4n0_49));
adder_full fa390(.sum(ws1b2n0_50), .c_out(ws1b2n1_49), .a(ws0b3n0_50), .b(ws0b3n1_50), .c_in(ws0b4n0_50));
adder_full fa391(.sum(ws1b2n0_51), .c_out(ws1b2n1_50), .a(ws0b3n0_51), .b(ws0b3n1_51), .c_in(ws0b4n0_51));
adder_half ha25(.sum(ws1b2n0_52), .c_out(ws1b2n1_51), .a(ws0b3n0_52), .b(ws0b3n1_52));
assign ws1b2n0_53 = ws0b3n0_53;
assign ws1b2n0_54 = ws0b3n0_54;
adder_half ha26(.sum(ws1b3n0_15), .c_out(ws1b3n1_14), .a(ws0b5n0_15), .b(ws0b5n1_15));
adder_half ha27(.sum(ws1b3n0_16), .c_out(ws1b3n1_15), .a(ws0b5n0_16), .b(ws0b5n1_16));
adder_half ha28(.sum(ws1b3n0_17), .c_out(ws1b3n1_16), .a(ws0b5n0_17), .b(ws0b5n1_17));
adder_full fa392(.sum(ws1b3n0_18), .c_out(ws1b3n1_17), .a(ws0b4n1_18), .b(ws0b5n0_18), .c_in(ws0b5n1_18));
adder_full fa393(.sum(ws1b3n0_19), .c_out(ws1b3n1_18), .a(ws0b4n1_19), .b(ws0b5n0_19), .c_in(ws0b5n1_19));
adder_full fa394(.sum(ws1b3n0_20), .c_out(ws1b3n1_19), .a(ws0b4n1_20), .b(ws0b5n0_20), .c_in(ws0b5n1_20));
adder_full fa395(.sum(ws1b3n0_21), .c_out(ws1b3n1_20), .a(ws0b4n1_21), .b(ws0b5n0_21), .c_in(ws0b5n1_21));
adder_full fa396(.sum(ws1b3n0_22), .c_out(ws1b3n1_21), .a(ws0b4n1_22), .b(ws0b5n0_22), .c_in(ws0b5n1_22));
adder_full fa397(.sum(ws1b3n0_23), .c_out(ws1b3n1_22), .a(ws0b4n1_23), .b(ws0b5n0_23), .c_in(ws0b5n1_23));
adder_full fa398(.sum(ws1b3n0_24), .c_out(ws1b3n1_23), .a(ws0b4n1_24), .b(ws0b5n0_24), .c_in(ws0b5n1_24));
adder_full fa399(.sum(ws1b3n0_25), .c_out(ws1b3n1_24), .a(ws0b4n1_25), .b(ws0b5n0_25), .c_in(ws0b5n1_25));
adder_full fa400(.sum(ws1b3n0_26), .c_out(ws1b3n1_25), .a(ws0b4n1_26), .b(ws0b5n0_26), .c_in(ws0b5n1_26));
adder_full fa401(.sum(ws1b3n0_27), .c_out(ws1b3n1_26), .a(ws0b4n1_27), .b(ws0b5n0_27), .c_in(ws0b5n1_27));
adder_full fa402(.sum(ws1b3n0_28), .c_out(ws1b3n1_27), .a(ws0b4n1_28), .b(ws0b5n0_28), .c_in(ws0b5n1_28));
adder_full fa403(.sum(ws1b3n0_29), .c_out(ws1b3n1_28), .a(ws0b4n1_29), .b(ws0b5n0_29), .c_in(ws0b5n1_29));
adder_full fa404(.sum(ws1b3n0_30), .c_out(ws1b3n1_29), .a(ws0b4n1_30), .b(ws0b5n0_30), .c_in(ws0b5n1_30));
adder_full fa405(.sum(ws1b3n0_31), .c_out(ws1b3n1_30), .a(ws0b4n1_31), .b(ws0b5n0_31), .c_in(ws0b5n1_31));
adder_full fa406(.sum(ws1b3n0_32), .c_out(ws1b3n1_31), .a(ws0b4n1_32), .b(ws0b5n0_32), .c_in(ws0b5n1_32));
adder_full fa407(.sum(ws1b3n0_33), .c_out(ws1b3n1_32), .a(ws0b4n1_33), .b(ws0b5n0_33), .c_in(ws0b5n1_33));
adder_full fa408(.sum(ws1b3n0_34), .c_out(ws1b3n1_33), .a(ws0b4n1_34), .b(ws0b5n0_34), .c_in(ws0b5n1_34));
adder_full fa409(.sum(ws1b3n0_35), .c_out(ws1b3n1_34), .a(ws0b4n1_35), .b(ws0b5n0_35), .c_in(ws0b5n1_35));
adder_full fa410(.sum(ws1b3n0_36), .c_out(ws1b3n1_35), .a(ws0b4n1_36), .b(ws0b5n0_36), .c_in(ws0b5n1_36));
adder_full fa411(.sum(ws1b3n0_37), .c_out(ws1b3n1_36), .a(ws0b4n1_37), .b(ws0b5n0_37), .c_in(ws0b5n1_37));
adder_full fa412(.sum(ws1b3n0_38), .c_out(ws1b3n1_37), .a(ws0b4n1_38), .b(ws0b5n0_38), .c_in(ws0b5n1_38));
adder_full fa413(.sum(ws1b3n0_39), .c_out(ws1b3n1_38), .a(ws0b4n1_39), .b(ws0b5n0_39), .c_in(ws0b5n1_39));
adder_full fa414(.sum(ws1b3n0_40), .c_out(ws1b3n1_39), .a(ws0b4n1_40), .b(ws0b5n0_40), .c_in(ws0b5n1_40));
adder_full fa415(.sum(ws1b3n0_41), .c_out(ws1b3n1_40), .a(ws0b4n1_41), .b(ws0b5n0_41), .c_in(ws0b5n1_41));
adder_full fa416(.sum(ws1b3n0_42), .c_out(ws1b3n1_41), .a(ws0b4n1_42), .b(ws0b5n0_42), .c_in(ws0b5n1_42));
adder_full fa417(.sum(ws1b3n0_43), .c_out(ws1b3n1_42), .a(ws0b4n1_43), .b(ws0b5n0_43), .c_in(ws0b5n1_43));
adder_full fa418(.sum(ws1b3n0_44), .c_out(ws1b3n1_43), .a(ws0b4n1_44), .b(ws0b5n0_44), .c_in(ws0b5n1_44));
adder_full fa419(.sum(ws1b3n0_45), .c_out(ws1b3n1_44), .a(ws0b4n1_45), .b(ws0b5n0_45), .c_in(ws0b5n1_45));
adder_full fa420(.sum(ws1b3n0_46), .c_out(ws1b3n1_45), .a(ws0b4n1_46), .b(ws0b5n0_46), .c_in(ws0b5n1_46));
adder_half ha29(.sum(ws1b3n0_47), .c_out(ws1b3n1_46), .a(ws0b4n1_47), .b(ws0b5n0_47));
adder_half ha30(.sum(ws1b3n0_48), .c_out(ws1b3n1_47), .a(ws0b4n1_48), .b(ws0b5n0_48));
assign ws1b3n0_49 = ws0b4n1_49;
assign ws1b4n0_9 = ws0b7n0_9;
assign ws1b4n0_10 = ws0b7n0_10;
assign ws1b4n0_11 = ws0b7n0_11;
adder_full fa421(.sum(ws1b4n0_12), .c_out(ws1b4n1_11), .a(ws0b6n0_12), .b(ws0b6n1_12), .c_in(ws0b7n0_12));
adder_full fa422(.sum(ws1b4n0_13), .c_out(ws1b4n1_12), .a(ws0b6n0_13), .b(ws0b6n1_13), .c_in(ws0b7n0_13));
adder_full fa423(.sum(ws1b4n0_14), .c_out(ws1b4n1_13), .a(ws0b6n0_14), .b(ws0b6n1_14), .c_in(ws0b7n0_14));
adder_full fa424(.sum(ws1b4n0_15), .c_out(ws1b4n1_14), .a(ws0b6n0_15), .b(ws0b6n1_15), .c_in(ws0b7n0_15));
adder_full fa425(.sum(ws1b4n0_16), .c_out(ws1b4n1_15), .a(ws0b6n0_16), .b(ws0b6n1_16), .c_in(ws0b7n0_16));
adder_full fa426(.sum(ws1b4n0_17), .c_out(ws1b4n1_16), .a(ws0b6n0_17), .b(ws0b6n1_17), .c_in(ws0b7n0_17));
adder_full fa427(.sum(ws1b4n0_18), .c_out(ws1b4n1_17), .a(ws0b6n0_18), .b(ws0b6n1_18), .c_in(ws0b7n0_18));
adder_full fa428(.sum(ws1b4n0_19), .c_out(ws1b4n1_18), .a(ws0b6n0_19), .b(ws0b6n1_19), .c_in(ws0b7n0_19));
adder_full fa429(.sum(ws1b4n0_20), .c_out(ws1b4n1_19), .a(ws0b6n0_20), .b(ws0b6n1_20), .c_in(ws0b7n0_20));
adder_full fa430(.sum(ws1b4n0_21), .c_out(ws1b4n1_20), .a(ws0b6n0_21), .b(ws0b6n1_21), .c_in(ws0b7n0_21));
adder_full fa431(.sum(ws1b4n0_22), .c_out(ws1b4n1_21), .a(ws0b6n0_22), .b(ws0b6n1_22), .c_in(ws0b7n0_22));
adder_full fa432(.sum(ws1b4n0_23), .c_out(ws1b4n1_22), .a(ws0b6n0_23), .b(ws0b6n1_23), .c_in(ws0b7n0_23));
adder_full fa433(.sum(ws1b4n0_24), .c_out(ws1b4n1_23), .a(ws0b6n0_24), .b(ws0b6n1_24), .c_in(ws0b7n0_24));
adder_full fa434(.sum(ws1b4n0_25), .c_out(ws1b4n1_24), .a(ws0b6n0_25), .b(ws0b6n1_25), .c_in(ws0b7n0_25));
adder_full fa435(.sum(ws1b4n0_26), .c_out(ws1b4n1_25), .a(ws0b6n0_26), .b(ws0b6n1_26), .c_in(ws0b7n0_26));
adder_full fa436(.sum(ws1b4n0_27), .c_out(ws1b4n1_26), .a(ws0b6n0_27), .b(ws0b6n1_27), .c_in(ws0b7n0_27));
adder_full fa437(.sum(ws1b4n0_28), .c_out(ws1b4n1_27), .a(ws0b6n0_28), .b(ws0b6n1_28), .c_in(ws0b7n0_28));
adder_full fa438(.sum(ws1b4n0_29), .c_out(ws1b4n1_28), .a(ws0b6n0_29), .b(ws0b6n1_29), .c_in(ws0b7n0_29));
adder_full fa439(.sum(ws1b4n0_30), .c_out(ws1b4n1_29), .a(ws0b6n0_30), .b(ws0b6n1_30), .c_in(ws0b7n0_30));
adder_full fa440(.sum(ws1b4n0_31), .c_out(ws1b4n1_30), .a(ws0b6n0_31), .b(ws0b6n1_31), .c_in(ws0b7n0_31));
adder_full fa441(.sum(ws1b4n0_32), .c_out(ws1b4n1_31), .a(ws0b6n0_32), .b(ws0b6n1_32), .c_in(ws0b7n0_32));
adder_full fa442(.sum(ws1b4n0_33), .c_out(ws1b4n1_32), .a(ws0b6n0_33), .b(ws0b6n1_33), .c_in(ws0b7n0_33));
adder_full fa443(.sum(ws1b4n0_34), .c_out(ws1b4n1_33), .a(ws0b6n0_34), .b(ws0b6n1_34), .c_in(ws0b7n0_34));
adder_full fa444(.sum(ws1b4n0_35), .c_out(ws1b4n1_34), .a(ws0b6n0_35), .b(ws0b6n1_35), .c_in(ws0b7n0_35));
adder_full fa445(.sum(ws1b4n0_36), .c_out(ws1b4n1_35), .a(ws0b6n0_36), .b(ws0b6n1_36), .c_in(ws0b7n0_36));
adder_full fa446(.sum(ws1b4n0_37), .c_out(ws1b4n1_36), .a(ws0b6n0_37), .b(ws0b6n1_37), .c_in(ws0b7n0_37));
adder_full fa447(.sum(ws1b4n0_38), .c_out(ws1b4n1_37), .a(ws0b6n0_38), .b(ws0b6n1_38), .c_in(ws0b7n0_38));
adder_full fa448(.sum(ws1b4n0_39), .c_out(ws1b4n1_38), .a(ws0b6n0_39), .b(ws0b6n1_39), .c_in(ws0b7n0_39));
adder_full fa449(.sum(ws1b4n0_40), .c_out(ws1b4n1_39), .a(ws0b6n0_40), .b(ws0b6n1_40), .c_in(ws0b7n0_40));
adder_full fa450(.sum(ws1b4n0_41), .c_out(ws1b4n1_40), .a(ws0b6n0_41), .b(ws0b6n1_41), .c_in(ws0b7n0_41));
adder_full fa451(.sum(ws1b4n0_42), .c_out(ws1b4n1_41), .a(ws0b6n0_42), .b(ws0b6n1_42), .c_in(ws0b7n0_42));
adder_half ha31(.sum(ws1b4n0_43), .c_out(ws1b4n1_42), .a(ws0b6n0_43), .b(ws0b6n1_43));
assign ws1b4n0_44 = ws0b6n0_44;
assign ws1b4n0_45 = ws0b6n0_45;
adder_half ha32(.sum(ws1b5n0_6), .c_out(ws1b5n1_5), .a(ws0b8n0_6), .b(ws0b8n1_6));
adder_half ha33(.sum(ws1b5n0_7), .c_out(ws1b5n1_6), .a(ws0b8n0_7), .b(ws0b8n1_7));
adder_half ha34(.sum(ws1b5n0_8), .c_out(ws1b5n1_7), .a(ws0b8n0_8), .b(ws0b8n1_8));
adder_full fa452(.sum(ws1b5n0_9), .c_out(ws1b5n1_8), .a(ws0b7n1_9), .b(ws0b8n0_9), .c_in(ws0b8n1_9));
adder_full fa453(.sum(ws1b5n0_10), .c_out(ws1b5n1_9), .a(ws0b7n1_10), .b(ws0b8n0_10), .c_in(ws0b8n1_10));
adder_full fa454(.sum(ws1b5n0_11), .c_out(ws1b5n1_10), .a(ws0b7n1_11), .b(ws0b8n0_11), .c_in(ws0b8n1_11));
adder_full fa455(.sum(ws1b5n0_12), .c_out(ws1b5n1_11), .a(ws0b7n1_12), .b(ws0b8n0_12), .c_in(ws0b8n1_12));
adder_full fa456(.sum(ws1b5n0_13), .c_out(ws1b5n1_12), .a(ws0b7n1_13), .b(ws0b8n0_13), .c_in(ws0b8n1_13));
adder_full fa457(.sum(ws1b5n0_14), .c_out(ws1b5n1_13), .a(ws0b7n1_14), .b(ws0b8n0_14), .c_in(ws0b8n1_14));
adder_full fa458(.sum(ws1b5n0_15), .c_out(ws1b5n1_14), .a(ws0b7n1_15), .b(ws0b8n0_15), .c_in(ws0b8n1_15));
adder_full fa459(.sum(ws1b5n0_16), .c_out(ws1b5n1_15), .a(ws0b7n1_16), .b(ws0b8n0_16), .c_in(ws0b8n1_16));
adder_full fa460(.sum(ws1b5n0_17), .c_out(ws1b5n1_16), .a(ws0b7n1_17), .b(ws0b8n0_17), .c_in(ws0b8n1_17));
adder_full fa461(.sum(ws1b5n0_18), .c_out(ws1b5n1_17), .a(ws0b7n1_18), .b(ws0b8n0_18), .c_in(ws0b8n1_18));
adder_full fa462(.sum(ws1b5n0_19), .c_out(ws1b5n1_18), .a(ws0b7n1_19), .b(ws0b8n0_19), .c_in(ws0b8n1_19));
adder_full fa463(.sum(ws1b5n0_20), .c_out(ws1b5n1_19), .a(ws0b7n1_20), .b(ws0b8n0_20), .c_in(ws0b8n1_20));
adder_full fa464(.sum(ws1b5n0_21), .c_out(ws1b5n1_20), .a(ws0b7n1_21), .b(ws0b8n0_21), .c_in(ws0b8n1_21));
adder_full fa465(.sum(ws1b5n0_22), .c_out(ws1b5n1_21), .a(ws0b7n1_22), .b(ws0b8n0_22), .c_in(ws0b8n1_22));
adder_full fa466(.sum(ws1b5n0_23), .c_out(ws1b5n1_22), .a(ws0b7n1_23), .b(ws0b8n0_23), .c_in(ws0b8n1_23));
adder_full fa467(.sum(ws1b5n0_24), .c_out(ws1b5n1_23), .a(ws0b7n1_24), .b(ws0b8n0_24), .c_in(ws0b8n1_24));
adder_full fa468(.sum(ws1b5n0_25), .c_out(ws1b5n1_24), .a(ws0b7n1_25), .b(ws0b8n0_25), .c_in(ws0b8n1_25));
adder_full fa469(.sum(ws1b5n0_26), .c_out(ws1b5n1_25), .a(ws0b7n1_26), .b(ws0b8n0_26), .c_in(ws0b8n1_26));
adder_full fa470(.sum(ws1b5n0_27), .c_out(ws1b5n1_26), .a(ws0b7n1_27), .b(ws0b8n0_27), .c_in(ws0b8n1_27));
adder_full fa471(.sum(ws1b5n0_28), .c_out(ws1b5n1_27), .a(ws0b7n1_28), .b(ws0b8n0_28), .c_in(ws0b8n1_28));
adder_full fa472(.sum(ws1b5n0_29), .c_out(ws1b5n1_28), .a(ws0b7n1_29), .b(ws0b8n0_29), .c_in(ws0b8n1_29));
adder_full fa473(.sum(ws1b5n0_30), .c_out(ws1b5n1_29), .a(ws0b7n1_30), .b(ws0b8n0_30), .c_in(ws0b8n1_30));
adder_full fa474(.sum(ws1b5n0_31), .c_out(ws1b5n1_30), .a(ws0b7n1_31), .b(ws0b8n0_31), .c_in(ws0b8n1_31));
adder_full fa475(.sum(ws1b5n0_32), .c_out(ws1b5n1_31), .a(ws0b7n1_32), .b(ws0b8n0_32), .c_in(ws0b8n1_32));
adder_full fa476(.sum(ws1b5n0_33), .c_out(ws1b5n1_32), .a(ws0b7n1_33), .b(ws0b8n0_33), .c_in(ws0b8n1_33));
adder_full fa477(.sum(ws1b5n0_34), .c_out(ws1b5n1_33), .a(ws0b7n1_34), .b(ws0b8n0_34), .c_in(ws0b8n1_34));
adder_full fa478(.sum(ws1b5n0_35), .c_out(ws1b5n1_34), .a(ws0b7n1_35), .b(ws0b8n0_35), .c_in(ws0b8n1_35));
adder_full fa479(.sum(ws1b5n0_36), .c_out(ws1b5n1_35), .a(ws0b7n1_36), .b(ws0b8n0_36), .c_in(ws0b8n1_36));
adder_full fa480(.sum(ws1b5n0_37), .c_out(ws1b5n1_36), .a(ws0b7n1_37), .b(ws0b8n0_37), .c_in(ws0b8n1_37));
adder_half ha35(.sum(ws1b5n0_38), .c_out(ws1b5n1_37), .a(ws0b7n1_38), .b(ws0b8n0_38));
adder_half ha36(.sum(ws1b5n0_39), .c_out(ws1b5n1_38), .a(ws0b7n1_39), .b(ws0b8n0_39));
assign ws1b5n0_40 = ws0b7n1_40;
assign ws1b6n0_2 = wand31_30;
adder_full fa481(.sum(ws1b6n0_3), .c_out(ws1b6n1_2), .a(ws0b9n0_3), .b(ws0b9n1_3), .c_in(wand30_30));
adder_full fa482(.sum(ws1b6n0_4), .c_out(ws1b6n1_3), .a(ws0b9n0_4), .b(ws0b9n1_4), .c_in(wand29_30));
adder_full fa483(.sum(ws1b6n0_5), .c_out(ws1b6n1_4), .a(ws0b9n0_5), .b(ws0b9n1_5), .c_in(wand28_30));
adder_full fa484(.sum(ws1b6n0_6), .c_out(ws1b6n1_5), .a(ws0b9n0_6), .b(ws0b9n1_6), .c_in(wand27_30));
adder_full fa485(.sum(ws1b6n0_7), .c_out(ws1b6n1_6), .a(ws0b9n0_7), .b(ws0b9n1_7), .c_in(wand26_30));
adder_full fa486(.sum(ws1b6n0_8), .c_out(ws1b6n1_7), .a(ws0b9n0_8), .b(ws0b9n1_8), .c_in(wand25_30));
adder_full fa487(.sum(ws1b6n0_9), .c_out(ws1b6n1_8), .a(ws0b9n0_9), .b(ws0b9n1_9), .c_in(wand24_30));
adder_full fa488(.sum(ws1b6n0_10), .c_out(ws1b6n1_9), .a(ws0b9n0_10), .b(ws0b9n1_10), .c_in(wand23_30));
adder_full fa489(.sum(ws1b6n0_11), .c_out(ws1b6n1_10), .a(ws0b9n0_11), .b(ws0b9n1_11), .c_in(wand22_30));
adder_full fa490(.sum(ws1b6n0_12), .c_out(ws1b6n1_11), .a(ws0b9n0_12), .b(ws0b9n1_12), .c_in(wand21_30));
adder_full fa491(.sum(ws1b6n0_13), .c_out(ws1b6n1_12), .a(ws0b9n0_13), .b(ws0b9n1_13), .c_in(wand20_30));
adder_full fa492(.sum(ws1b6n0_14), .c_out(ws1b6n1_13), .a(ws0b9n0_14), .b(ws0b9n1_14), .c_in(wand19_30));
adder_full fa493(.sum(ws1b6n0_15), .c_out(ws1b6n1_14), .a(ws0b9n0_15), .b(ws0b9n1_15), .c_in(wand18_30));
adder_full fa494(.sum(ws1b6n0_16), .c_out(ws1b6n1_15), .a(ws0b9n0_16), .b(ws0b9n1_16), .c_in(wand17_30));
adder_full fa495(.sum(ws1b6n0_17), .c_out(ws1b6n1_16), .a(ws0b9n0_17), .b(ws0b9n1_17), .c_in(wand16_30));
adder_full fa496(.sum(ws1b6n0_18), .c_out(ws1b6n1_17), .a(ws0b9n0_18), .b(ws0b9n1_18), .c_in(wand15_30));
adder_full fa497(.sum(ws1b6n0_19), .c_out(ws1b6n1_18), .a(ws0b9n0_19), .b(ws0b9n1_19), .c_in(wand14_30));
adder_full fa498(.sum(ws1b6n0_20), .c_out(ws1b6n1_19), .a(ws0b9n0_20), .b(ws0b9n1_20), .c_in(wand13_30));
adder_full fa499(.sum(ws1b6n0_21), .c_out(ws1b6n1_20), .a(ws0b9n0_21), .b(ws0b9n1_21), .c_in(wand12_30));
adder_full fa500(.sum(ws1b6n0_22), .c_out(ws1b6n1_21), .a(ws0b9n0_22), .b(ws0b9n1_22), .c_in(wand11_30));
adder_full fa501(.sum(ws1b6n0_23), .c_out(ws1b6n1_22), .a(ws0b9n0_23), .b(ws0b9n1_23), .c_in(wand10_30));
adder_full fa502(.sum(ws1b6n0_24), .c_out(ws1b6n1_23), .a(ws0b9n0_24), .b(ws0b9n1_24), .c_in(wand9_30));
adder_full fa503(.sum(ws1b6n0_25), .c_out(ws1b6n1_24), .a(ws0b9n0_25), .b(ws0b9n1_25), .c_in(wand8_30));
adder_full fa504(.sum(ws1b6n0_26), .c_out(ws1b6n1_25), .a(ws0b9n0_26), .b(ws0b9n1_26), .c_in(wand7_30));
adder_full fa505(.sum(ws1b6n0_27), .c_out(ws1b6n1_26), .a(ws0b9n0_27), .b(ws0b9n1_27), .c_in(wand6_30));
adder_full fa506(.sum(ws1b6n0_28), .c_out(ws1b6n1_27), .a(ws0b9n0_28), .b(ws0b9n1_28), .c_in(wand5_30));
adder_full fa507(.sum(ws1b6n0_29), .c_out(ws1b6n1_28), .a(ws0b9n0_29), .b(ws0b9n1_29), .c_in(wand4_30));
adder_full fa508(.sum(ws1b6n0_30), .c_out(ws1b6n1_29), .a(ws0b9n0_30), .b(ws0b9n1_30), .c_in(wand3_30));
adder_full fa509(.sum(ws1b6n0_31), .c_out(ws1b6n1_30), .a(ws0b9n0_31), .b(ws0b9n1_31), .c_in(wand2_30));
adder_full fa510(.sum(ws1b6n0_32), .c_out(ws1b6n1_31), .a(ws0b9n0_32), .b(ws0b9n1_32), .c_in(wand1_30));
adder_full fa511(.sum(ws1b6n0_33), .c_out(ws1b6n1_32), .a(ws0b9n0_33), .b(ws0b9n1_33), .c_in(wand0_30));
adder_half ha37(.sum(ws1b6n0_34), .c_out(ws1b6n1_33), .a(ws0b9n0_34), .b(ws0b9n1_34));
assign ws1b6n0_35 = ws0b9n0_35;
assign ws1b6n0_36 = ws0b9n0_36;

assign ws2b0n0_24 = ws1b1n0_24;
assign ws2b0n0_25 = ws1b1n0_25;
assign ws2b0n0_26 = ws1b1n0_26;
adder_half ha38(.sum(ws2b0n0_27), .c_out(ws2b0n1_26), .a(ws1b0n0_27), .b(ws1b1n0_27));
adder_half ha39(.sum(ws2b0n0_28), .c_out(ws2b0n1_27), .a(ws1b0n0_28), .b(ws1b1n0_28));
adder_full fa512(.sum(ws2b0n0_29), .c_out(ws2b0n1_28), .a(ws1b0n0_29), .b(ws1b0n1_29), .c_in(ws1b1n0_29));
adder_full fa513(.sum(ws2b0n0_30), .c_out(ws2b0n1_29), .a(ws1b0n0_30), .b(ws1b0n1_30), .c_in(ws1b1n0_30));
adder_full fa514(.sum(ws2b0n0_31), .c_out(ws2b0n1_30), .a(ws1b0n0_31), .b(ws1b0n1_31), .c_in(ws1b1n0_31));
adder_full fa515(.sum(ws2b0n0_32), .c_out(ws2b0n1_31), .a(ws1b0n0_32), .b(ws1b0n1_32), .c_in(ws1b1n0_32));
adder_full fa516(.sum(ws2b0n0_33), .c_out(ws2b0n1_32), .a(ws1b0n0_33), .b(ws1b0n1_33), .c_in(ws1b1n0_33));
adder_full fa517(.sum(ws2b0n0_34), .c_out(ws2b0n1_33), .a(ws1b0n0_34), .b(ws1b0n1_34), .c_in(ws1b1n0_34));
adder_full fa518(.sum(ws2b0n0_35), .c_out(ws2b0n1_34), .a(ws1b0n0_35), .b(ws1b0n1_35), .c_in(ws1b1n0_35));
adder_full fa519(.sum(ws2b0n0_36), .c_out(ws2b0n1_35), .a(ws1b0n0_36), .b(ws1b0n1_36), .c_in(ws1b1n0_36));
adder_full fa520(.sum(ws2b0n0_37), .c_out(ws2b0n1_36), .a(ws1b0n0_37), .b(ws1b0n1_37), .c_in(ws1b1n0_37));
adder_full fa521(.sum(ws2b0n0_38), .c_out(ws2b0n1_37), .a(ws1b0n0_38), .b(ws1b0n1_38), .c_in(ws1b1n0_38));
adder_full fa522(.sum(ws2b0n0_39), .c_out(ws2b0n1_38), .a(ws1b0n0_39), .b(ws1b0n1_39), .c_in(ws1b1n0_39));
adder_full fa523(.sum(ws2b0n0_40), .c_out(ws2b0n1_39), .a(ws1b0n0_40), .b(ws1b0n1_40), .c_in(ws1b1n0_40));
adder_full fa524(.sum(ws2b0n0_41), .c_out(ws2b0n1_40), .a(ws1b0n0_41), .b(ws1b0n1_41), .c_in(ws1b1n0_41));
adder_full fa525(.sum(ws2b0n0_42), .c_out(ws2b0n1_41), .a(ws1b0n0_42), .b(ws1b0n1_42), .c_in(ws1b1n0_42));
adder_full fa526(.sum(ws2b0n0_43), .c_out(ws2b0n1_42), .a(ws1b0n0_43), .b(ws1b0n1_43), .c_in(ws1b1n0_43));
adder_full fa527(.sum(ws2b0n0_44), .c_out(ws2b0n1_43), .a(ws1b0n0_44), .b(ws1b0n1_44), .c_in(ws1b1n0_44));
adder_full fa528(.sum(ws2b0n0_45), .c_out(ws2b0n1_44), .a(ws1b0n0_45), .b(ws1b0n1_45), .c_in(ws1b1n0_45));
adder_full fa529(.sum(ws2b0n0_46), .c_out(ws2b0n1_45), .a(ws1b0n0_46), .b(ws1b0n1_46), .c_in(ws1b1n0_46));
adder_full fa530(.sum(ws2b0n0_47), .c_out(ws2b0n1_46), .a(ws1b0n0_47), .b(ws1b0n1_47), .c_in(ws1b1n0_47));
adder_full fa531(.sum(ws2b0n0_48), .c_out(ws2b0n1_47), .a(ws1b0n0_48), .b(ws1b0n1_48), .c_in(ws1b1n0_48));
adder_full fa532(.sum(ws2b0n0_49), .c_out(ws2b0n1_48), .a(ws1b0n0_49), .b(ws1b0n1_49), .c_in(ws1b1n0_49));
adder_full fa533(.sum(ws2b0n0_50), .c_out(ws2b0n1_49), .a(ws1b0n0_50), .b(ws1b0n1_50), .c_in(ws1b1n0_50));
adder_full fa534(.sum(ws2b0n0_51), .c_out(ws2b0n1_50), .a(ws1b0n0_51), .b(ws1b0n1_51), .c_in(ws1b1n0_51));
adder_full fa535(.sum(ws2b0n0_52), .c_out(ws2b0n1_51), .a(ws1b0n0_52), .b(ws1b0n1_52), .c_in(ws1b1n0_52));
adder_full fa536(.sum(ws2b0n0_53), .c_out(ws2b0n1_52), .a(ws1b0n0_53), .b(ws1b0n1_53), .c_in(ws1b1n0_53));
adder_full fa537(.sum(ws2b0n0_54), .c_out(ws2b0n1_53), .a(ws1b0n0_54), .b(ws1b0n1_54), .c_in(ws1b1n0_54));
adder_full fa538(.sum(ws2b0n0_55), .c_out(ws2b0n1_54), .a(ws1b0n0_55), .b(ws1b0n1_55), .c_in(ws1b1n0_55));
adder_full fa539(.sum(ws2b0n0_56), .c_out(ws2b0n1_55), .a(ws1b0n0_56), .b(ws1b0n1_56), .c_in(ws1b1n0_56));
adder_full fa540(.sum(ws2b0n0_57), .c_out(ws2b0n1_56), .a(ws1b0n0_57), .b(ws1b0n1_57), .c_in(ws1b1n0_57));
adder_full fa541(.sum(ws2b0n0_58), .c_out(ws2b0n1_57), .a(ws1b0n0_58), .b(ws1b0n1_58), .c_in(ws1b1n0_58));
adder_half ha40(.sum(ws2b0n0_59), .c_out(ws2b0n1_58), .a(ws1b0n0_59), .b(ws1b0n1_59));
adder_half ha41(.sum(ws2b0n0_60), .c_out(ws2b0n1_59), .a(ws1b0n0_60), .b(ws1b0n1_60));
assign ws2b0n0_61 = ws1b0n0_61;
assign ws2b0n0_62 = ws1b0n0_62;
assign ws2b0n0_63 = ws1b0n0_63;
assign ws2b1n0_18 = ws1b2n0_18;
assign ws2b1n0_19 = ws1b2n0_19;
adder_half ha42(.sum(ws2b1n0_20), .c_out(ws2b1n1_19), .a(ws1b2n0_20), .b(ws1b2n1_20));
adder_half ha43(.sum(ws2b1n0_21), .c_out(ws2b1n1_20), .a(ws1b2n0_21), .b(ws1b2n1_21));
adder_half ha44(.sum(ws2b1n0_22), .c_out(ws2b1n1_21), .a(ws1b2n0_22), .b(ws1b2n1_22));
adder_full fa542(.sum(ws2b1n0_23), .c_out(ws2b1n1_22), .a(ws1b1n1_23), .b(ws1b2n0_23), .c_in(ws1b2n1_23));
adder_full fa543(.sum(ws2b1n0_24), .c_out(ws2b1n1_23), .a(ws1b1n1_24), .b(ws1b2n0_24), .c_in(ws1b2n1_24));
adder_full fa544(.sum(ws2b1n0_25), .c_out(ws2b1n1_24), .a(ws1b1n1_25), .b(ws1b2n0_25), .c_in(ws1b2n1_25));
adder_full fa545(.sum(ws2b1n0_26), .c_out(ws2b1n1_25), .a(ws1b1n1_26), .b(ws1b2n0_26), .c_in(ws1b2n1_26));
adder_full fa546(.sum(ws2b1n0_27), .c_out(ws2b1n1_26), .a(ws1b1n1_27), .b(ws1b2n0_27), .c_in(ws1b2n1_27));
adder_full fa547(.sum(ws2b1n0_28), .c_out(ws2b1n1_27), .a(ws1b1n1_28), .b(ws1b2n0_28), .c_in(ws1b2n1_28));
adder_full fa548(.sum(ws2b1n0_29), .c_out(ws2b1n1_28), .a(ws1b1n1_29), .b(ws1b2n0_29), .c_in(ws1b2n1_29));
adder_full fa549(.sum(ws2b1n0_30), .c_out(ws2b1n1_29), .a(ws1b1n1_30), .b(ws1b2n0_30), .c_in(ws1b2n1_30));
adder_full fa550(.sum(ws2b1n0_31), .c_out(ws2b1n1_30), .a(ws1b1n1_31), .b(ws1b2n0_31), .c_in(ws1b2n1_31));
adder_full fa551(.sum(ws2b1n0_32), .c_out(ws2b1n1_31), .a(ws1b1n1_32), .b(ws1b2n0_32), .c_in(ws1b2n1_32));
adder_full fa552(.sum(ws2b1n0_33), .c_out(ws2b1n1_32), .a(ws1b1n1_33), .b(ws1b2n0_33), .c_in(ws1b2n1_33));
adder_full fa553(.sum(ws2b1n0_34), .c_out(ws2b1n1_33), .a(ws1b1n1_34), .b(ws1b2n0_34), .c_in(ws1b2n1_34));
adder_full fa554(.sum(ws2b1n0_35), .c_out(ws2b1n1_34), .a(ws1b1n1_35), .b(ws1b2n0_35), .c_in(ws1b2n1_35));
adder_full fa555(.sum(ws2b1n0_36), .c_out(ws2b1n1_35), .a(ws1b1n1_36), .b(ws1b2n0_36), .c_in(ws1b2n1_36));
adder_full fa556(.sum(ws2b1n0_37), .c_out(ws2b1n1_36), .a(ws1b1n1_37), .b(ws1b2n0_37), .c_in(ws1b2n1_37));
adder_full fa557(.sum(ws2b1n0_38), .c_out(ws2b1n1_37), .a(ws1b1n1_38), .b(ws1b2n0_38), .c_in(ws1b2n1_38));
adder_full fa558(.sum(ws2b1n0_39), .c_out(ws2b1n1_38), .a(ws1b1n1_39), .b(ws1b2n0_39), .c_in(ws1b2n1_39));
adder_full fa559(.sum(ws2b1n0_40), .c_out(ws2b1n1_39), .a(ws1b1n1_40), .b(ws1b2n0_40), .c_in(ws1b2n1_40));
adder_full fa560(.sum(ws2b1n0_41), .c_out(ws2b1n1_40), .a(ws1b1n1_41), .b(ws1b2n0_41), .c_in(ws1b2n1_41));
adder_full fa561(.sum(ws2b1n0_42), .c_out(ws2b1n1_41), .a(ws1b1n1_42), .b(ws1b2n0_42), .c_in(ws1b2n1_42));
adder_full fa562(.sum(ws2b1n0_43), .c_out(ws2b1n1_42), .a(ws1b1n1_43), .b(ws1b2n0_43), .c_in(ws1b2n1_43));
adder_full fa563(.sum(ws2b1n0_44), .c_out(ws2b1n1_43), .a(ws1b1n1_44), .b(ws1b2n0_44), .c_in(ws1b2n1_44));
adder_full fa564(.sum(ws2b1n0_45), .c_out(ws2b1n1_44), .a(ws1b1n1_45), .b(ws1b2n0_45), .c_in(ws1b2n1_45));
adder_full fa565(.sum(ws2b1n0_46), .c_out(ws2b1n1_45), .a(ws1b1n1_46), .b(ws1b2n0_46), .c_in(ws1b2n1_46));
adder_full fa566(.sum(ws2b1n0_47), .c_out(ws2b1n1_46), .a(ws1b1n1_47), .b(ws1b2n0_47), .c_in(ws1b2n1_47));
adder_full fa567(.sum(ws2b1n0_48), .c_out(ws2b1n1_47), .a(ws1b1n1_48), .b(ws1b2n0_48), .c_in(ws1b2n1_48));
adder_full fa568(.sum(ws2b1n0_49), .c_out(ws2b1n1_48), .a(ws1b1n1_49), .b(ws1b2n0_49), .c_in(ws1b2n1_49));
adder_full fa569(.sum(ws2b1n0_50), .c_out(ws2b1n1_49), .a(ws1b1n1_50), .b(ws1b2n0_50), .c_in(ws1b2n1_50));
adder_full fa570(.sum(ws2b1n0_51), .c_out(ws2b1n1_50), .a(ws1b1n1_51), .b(ws1b2n0_51), .c_in(ws1b2n1_51));
adder_half ha45(.sum(ws2b1n0_52), .c_out(ws2b1n1_51), .a(ws1b1n1_52), .b(ws1b2n0_52));
adder_half ha46(.sum(ws2b1n0_53), .c_out(ws2b1n1_52), .a(ws1b1n1_53), .b(ws1b2n0_53));
adder_half ha47(.sum(ws2b1n0_54), .c_out(ws2b1n1_53), .a(ws1b1n1_54), .b(ws1b2n0_54));
assign ws2b1n0_55 = ws1b1n1_55;
assign ws2b1n0_56 = ws1b1n1_56;
assign ws2b2n0_9 = ws1b4n0_9;
assign ws2b2n0_10 = ws1b4n0_10;
assign ws2b2n0_11 = ws1b4n0_11;
assign ws2b2n0_12 = ws1b4n0_12;
assign ws2b2n0_13 = ws1b4n0_13;
adder_half ha48(.sum(ws2b2n0_14), .c_out(ws2b2n1_13), .a(ws1b3n1_14), .b(ws1b4n0_14));
adder_full fa571(.sum(ws2b2n0_15), .c_out(ws2b2n1_14), .a(ws1b3n0_15), .b(ws1b3n1_15), .c_in(ws1b4n0_15));
adder_full fa572(.sum(ws2b2n0_16), .c_out(ws2b2n1_15), .a(ws1b3n0_16), .b(ws1b3n1_16), .c_in(ws1b4n0_16));
adder_full fa573(.sum(ws2b2n0_17), .c_out(ws2b2n1_16), .a(ws1b3n0_17), .b(ws1b3n1_17), .c_in(ws1b4n0_17));
adder_full fa574(.sum(ws2b2n0_18), .c_out(ws2b2n1_17), .a(ws1b3n0_18), .b(ws1b3n1_18), .c_in(ws1b4n0_18));
adder_full fa575(.sum(ws2b2n0_19), .c_out(ws2b2n1_18), .a(ws1b3n0_19), .b(ws1b3n1_19), .c_in(ws1b4n0_19));
adder_full fa576(.sum(ws2b2n0_20), .c_out(ws2b2n1_19), .a(ws1b3n0_20), .b(ws1b3n1_20), .c_in(ws1b4n0_20));
adder_full fa577(.sum(ws2b2n0_21), .c_out(ws2b2n1_20), .a(ws1b3n0_21), .b(ws1b3n1_21), .c_in(ws1b4n0_21));
adder_full fa578(.sum(ws2b2n0_22), .c_out(ws2b2n1_21), .a(ws1b3n0_22), .b(ws1b3n1_22), .c_in(ws1b4n0_22));
adder_full fa579(.sum(ws2b2n0_23), .c_out(ws2b2n1_22), .a(ws1b3n0_23), .b(ws1b3n1_23), .c_in(ws1b4n0_23));
adder_full fa580(.sum(ws2b2n0_24), .c_out(ws2b2n1_23), .a(ws1b3n0_24), .b(ws1b3n1_24), .c_in(ws1b4n0_24));
adder_full fa581(.sum(ws2b2n0_25), .c_out(ws2b2n1_24), .a(ws1b3n0_25), .b(ws1b3n1_25), .c_in(ws1b4n0_25));
adder_full fa582(.sum(ws2b2n0_26), .c_out(ws2b2n1_25), .a(ws1b3n0_26), .b(ws1b3n1_26), .c_in(ws1b4n0_26));
adder_full fa583(.sum(ws2b2n0_27), .c_out(ws2b2n1_26), .a(ws1b3n0_27), .b(ws1b3n1_27), .c_in(ws1b4n0_27));
adder_full fa584(.sum(ws2b2n0_28), .c_out(ws2b2n1_27), .a(ws1b3n0_28), .b(ws1b3n1_28), .c_in(ws1b4n0_28));
adder_full fa585(.sum(ws2b2n0_29), .c_out(ws2b2n1_28), .a(ws1b3n0_29), .b(ws1b3n1_29), .c_in(ws1b4n0_29));
adder_full fa586(.sum(ws2b2n0_30), .c_out(ws2b2n1_29), .a(ws1b3n0_30), .b(ws1b3n1_30), .c_in(ws1b4n0_30));
adder_full fa587(.sum(ws2b2n0_31), .c_out(ws2b2n1_30), .a(ws1b3n0_31), .b(ws1b3n1_31), .c_in(ws1b4n0_31));
adder_full fa588(.sum(ws2b2n0_32), .c_out(ws2b2n1_31), .a(ws1b3n0_32), .b(ws1b3n1_32), .c_in(ws1b4n0_32));
adder_full fa589(.sum(ws2b2n0_33), .c_out(ws2b2n1_32), .a(ws1b3n0_33), .b(ws1b3n1_33), .c_in(ws1b4n0_33));
adder_full fa590(.sum(ws2b2n0_34), .c_out(ws2b2n1_33), .a(ws1b3n0_34), .b(ws1b3n1_34), .c_in(ws1b4n0_34));
adder_full fa591(.sum(ws2b2n0_35), .c_out(ws2b2n1_34), .a(ws1b3n0_35), .b(ws1b3n1_35), .c_in(ws1b4n0_35));
adder_full fa592(.sum(ws2b2n0_36), .c_out(ws2b2n1_35), .a(ws1b3n0_36), .b(ws1b3n1_36), .c_in(ws1b4n0_36));
adder_full fa593(.sum(ws2b2n0_37), .c_out(ws2b2n1_36), .a(ws1b3n0_37), .b(ws1b3n1_37), .c_in(ws1b4n0_37));
adder_full fa594(.sum(ws2b2n0_38), .c_out(ws2b2n1_37), .a(ws1b3n0_38), .b(ws1b3n1_38), .c_in(ws1b4n0_38));
adder_full fa595(.sum(ws2b2n0_39), .c_out(ws2b2n1_38), .a(ws1b3n0_39), .b(ws1b3n1_39), .c_in(ws1b4n0_39));
adder_full fa596(.sum(ws2b2n0_40), .c_out(ws2b2n1_39), .a(ws1b3n0_40), .b(ws1b3n1_40), .c_in(ws1b4n0_40));
adder_full fa597(.sum(ws2b2n0_41), .c_out(ws2b2n1_40), .a(ws1b3n0_41), .b(ws1b3n1_41), .c_in(ws1b4n0_41));
adder_full fa598(.sum(ws2b2n0_42), .c_out(ws2b2n1_41), .a(ws1b3n0_42), .b(ws1b3n1_42), .c_in(ws1b4n0_42));
adder_full fa599(.sum(ws2b2n0_43), .c_out(ws2b2n1_42), .a(ws1b3n0_43), .b(ws1b3n1_43), .c_in(ws1b4n0_43));
adder_full fa600(.sum(ws2b2n0_44), .c_out(ws2b2n1_43), .a(ws1b3n0_44), .b(ws1b3n1_44), .c_in(ws1b4n0_44));
adder_full fa601(.sum(ws2b2n0_45), .c_out(ws2b2n1_44), .a(ws1b3n0_45), .b(ws1b3n1_45), .c_in(ws1b4n0_45));
adder_half ha49(.sum(ws2b2n0_46), .c_out(ws2b2n1_45), .a(ws1b3n0_46), .b(ws1b3n1_46));
adder_half ha50(.sum(ws2b2n0_47), .c_out(ws2b2n1_46), .a(ws1b3n0_47), .b(ws1b3n1_47));
assign ws2b2n0_48 = ws1b3n0_48;
assign ws2b2n0_49 = ws1b3n0_49;
assign ws2b3n0_5 = ws1b5n1_5;
adder_half ha51(.sum(ws2b3n0_6), .c_out(ws2b3n1_5), .a(ws1b5n0_6), .b(ws1b5n1_6));
adder_half ha52(.sum(ws2b3n0_7), .c_out(ws2b3n1_6), .a(ws1b5n0_7), .b(ws1b5n1_7));
adder_half ha53(.sum(ws2b3n0_8), .c_out(ws2b3n1_7), .a(ws1b5n0_8), .b(ws1b5n1_8));
adder_half ha54(.sum(ws2b3n0_9), .c_out(ws2b3n1_8), .a(ws1b5n0_9), .b(ws1b5n1_9));
adder_half ha55(.sum(ws2b3n0_10), .c_out(ws2b3n1_9), .a(ws1b5n0_10), .b(ws1b5n1_10));
adder_full fa602(.sum(ws2b3n0_11), .c_out(ws2b3n1_10), .a(ws1b4n1_11), .b(ws1b5n0_11), .c_in(ws1b5n1_11));
adder_full fa603(.sum(ws2b3n0_12), .c_out(ws2b3n1_11), .a(ws1b4n1_12), .b(ws1b5n0_12), .c_in(ws1b5n1_12));
adder_full fa604(.sum(ws2b3n0_13), .c_out(ws2b3n1_12), .a(ws1b4n1_13), .b(ws1b5n0_13), .c_in(ws1b5n1_13));
adder_full fa605(.sum(ws2b3n0_14), .c_out(ws2b3n1_13), .a(ws1b4n1_14), .b(ws1b5n0_14), .c_in(ws1b5n1_14));
adder_full fa606(.sum(ws2b3n0_15), .c_out(ws2b3n1_14), .a(ws1b4n1_15), .b(ws1b5n0_15), .c_in(ws1b5n1_15));
adder_full fa607(.sum(ws2b3n0_16), .c_out(ws2b3n1_15), .a(ws1b4n1_16), .b(ws1b5n0_16), .c_in(ws1b5n1_16));
adder_full fa608(.sum(ws2b3n0_17), .c_out(ws2b3n1_16), .a(ws1b4n1_17), .b(ws1b5n0_17), .c_in(ws1b5n1_17));
adder_full fa609(.sum(ws2b3n0_18), .c_out(ws2b3n1_17), .a(ws1b4n1_18), .b(ws1b5n0_18), .c_in(ws1b5n1_18));
adder_full fa610(.sum(ws2b3n0_19), .c_out(ws2b3n1_18), .a(ws1b4n1_19), .b(ws1b5n0_19), .c_in(ws1b5n1_19));
adder_full fa611(.sum(ws2b3n0_20), .c_out(ws2b3n1_19), .a(ws1b4n1_20), .b(ws1b5n0_20), .c_in(ws1b5n1_20));
adder_full fa612(.sum(ws2b3n0_21), .c_out(ws2b3n1_20), .a(ws1b4n1_21), .b(ws1b5n0_21), .c_in(ws1b5n1_21));
adder_full fa613(.sum(ws2b3n0_22), .c_out(ws2b3n1_21), .a(ws1b4n1_22), .b(ws1b5n0_22), .c_in(ws1b5n1_22));
adder_full fa614(.sum(ws2b3n0_23), .c_out(ws2b3n1_22), .a(ws1b4n1_23), .b(ws1b5n0_23), .c_in(ws1b5n1_23));
adder_full fa615(.sum(ws2b3n0_24), .c_out(ws2b3n1_23), .a(ws1b4n1_24), .b(ws1b5n0_24), .c_in(ws1b5n1_24));
adder_full fa616(.sum(ws2b3n0_25), .c_out(ws2b3n1_24), .a(ws1b4n1_25), .b(ws1b5n0_25), .c_in(ws1b5n1_25));
adder_full fa617(.sum(ws2b3n0_26), .c_out(ws2b3n1_25), .a(ws1b4n1_26), .b(ws1b5n0_26), .c_in(ws1b5n1_26));
adder_full fa618(.sum(ws2b3n0_27), .c_out(ws2b3n1_26), .a(ws1b4n1_27), .b(ws1b5n0_27), .c_in(ws1b5n1_27));
adder_full fa619(.sum(ws2b3n0_28), .c_out(ws2b3n1_27), .a(ws1b4n1_28), .b(ws1b5n0_28), .c_in(ws1b5n1_28));
adder_full fa620(.sum(ws2b3n0_29), .c_out(ws2b3n1_28), .a(ws1b4n1_29), .b(ws1b5n0_29), .c_in(ws1b5n1_29));
adder_full fa621(.sum(ws2b3n0_30), .c_out(ws2b3n1_29), .a(ws1b4n1_30), .b(ws1b5n0_30), .c_in(ws1b5n1_30));
adder_full fa622(.sum(ws2b3n0_31), .c_out(ws2b3n1_30), .a(ws1b4n1_31), .b(ws1b5n0_31), .c_in(ws1b5n1_31));
adder_full fa623(.sum(ws2b3n0_32), .c_out(ws2b3n1_31), .a(ws1b4n1_32), .b(ws1b5n0_32), .c_in(ws1b5n1_32));
adder_full fa624(.sum(ws2b3n0_33), .c_out(ws2b3n1_32), .a(ws1b4n1_33), .b(ws1b5n0_33), .c_in(ws1b5n1_33));
adder_full fa625(.sum(ws2b3n0_34), .c_out(ws2b3n1_33), .a(ws1b4n1_34), .b(ws1b5n0_34), .c_in(ws1b5n1_34));
adder_full fa626(.sum(ws2b3n0_35), .c_out(ws2b3n1_34), .a(ws1b4n1_35), .b(ws1b5n0_35), .c_in(ws1b5n1_35));
adder_full fa627(.sum(ws2b3n0_36), .c_out(ws2b3n1_35), .a(ws1b4n1_36), .b(ws1b5n0_36), .c_in(ws1b5n1_36));
adder_full fa628(.sum(ws2b3n0_37), .c_out(ws2b3n1_36), .a(ws1b4n1_37), .b(ws1b5n0_37), .c_in(ws1b5n1_37));
adder_full fa629(.sum(ws2b3n0_38), .c_out(ws2b3n1_37), .a(ws1b4n1_38), .b(ws1b5n0_38), .c_in(ws1b5n1_38));
adder_half ha56(.sum(ws2b3n0_39), .c_out(ws2b3n1_38), .a(ws1b4n1_39), .b(ws1b5n0_39));
adder_half ha57(.sum(ws2b3n0_40), .c_out(ws2b3n1_39), .a(ws1b4n1_40), .b(ws1b5n0_40));
assign ws2b3n0_41 = ws1b4n1_41;
assign ws2b3n0_42 = ws1b4n1_42;
assign ws2b4n0_1 = wand31_31;
adder_full fa630(.sum(ws2b4n0_2), .c_out(ws2b4n1_1), .a(ws1b6n0_2), .b(ws1b6n1_2), .c_in(wand30_31));
adder_full fa631(.sum(ws2b4n0_3), .c_out(ws2b4n1_2), .a(ws1b6n0_3), .b(ws1b6n1_3), .c_in(wand29_31));
adder_full fa632(.sum(ws2b4n0_4), .c_out(ws2b4n1_3), .a(ws1b6n0_4), .b(ws1b6n1_4), .c_in(wand28_31));
adder_full fa633(.sum(ws2b4n0_5), .c_out(ws2b4n1_4), .a(ws1b6n0_5), .b(ws1b6n1_5), .c_in(wand27_31));
adder_full fa634(.sum(ws2b4n0_6), .c_out(ws2b4n1_5), .a(ws1b6n0_6), .b(ws1b6n1_6), .c_in(wand26_31));
adder_full fa635(.sum(ws2b4n0_7), .c_out(ws2b4n1_6), .a(ws1b6n0_7), .b(ws1b6n1_7), .c_in(wand25_31));
adder_full fa636(.sum(ws2b4n0_8), .c_out(ws2b4n1_7), .a(ws1b6n0_8), .b(ws1b6n1_8), .c_in(wand24_31));
adder_full fa637(.sum(ws2b4n0_9), .c_out(ws2b4n1_8), .a(ws1b6n0_9), .b(ws1b6n1_9), .c_in(wand23_31));
adder_full fa638(.sum(ws2b4n0_10), .c_out(ws2b4n1_9), .a(ws1b6n0_10), .b(ws1b6n1_10), .c_in(wand22_31));
adder_full fa639(.sum(ws2b4n0_11), .c_out(ws2b4n1_10), .a(ws1b6n0_11), .b(ws1b6n1_11), .c_in(wand21_31));
adder_full fa640(.sum(ws2b4n0_12), .c_out(ws2b4n1_11), .a(ws1b6n0_12), .b(ws1b6n1_12), .c_in(wand20_31));
adder_full fa641(.sum(ws2b4n0_13), .c_out(ws2b4n1_12), .a(ws1b6n0_13), .b(ws1b6n1_13), .c_in(wand19_31));
adder_full fa642(.sum(ws2b4n0_14), .c_out(ws2b4n1_13), .a(ws1b6n0_14), .b(ws1b6n1_14), .c_in(wand18_31));
adder_full fa643(.sum(ws2b4n0_15), .c_out(ws2b4n1_14), .a(ws1b6n0_15), .b(ws1b6n1_15), .c_in(wand17_31));
adder_full fa644(.sum(ws2b4n0_16), .c_out(ws2b4n1_15), .a(ws1b6n0_16), .b(ws1b6n1_16), .c_in(wand16_31));
adder_full fa645(.sum(ws2b4n0_17), .c_out(ws2b4n1_16), .a(ws1b6n0_17), .b(ws1b6n1_17), .c_in(wand15_31));
adder_full fa646(.sum(ws2b4n0_18), .c_out(ws2b4n1_17), .a(ws1b6n0_18), .b(ws1b6n1_18), .c_in(wand14_31));
adder_full fa647(.sum(ws2b4n0_19), .c_out(ws2b4n1_18), .a(ws1b6n0_19), .b(ws1b6n1_19), .c_in(wand13_31));
adder_full fa648(.sum(ws2b4n0_20), .c_out(ws2b4n1_19), .a(ws1b6n0_20), .b(ws1b6n1_20), .c_in(wand12_31));
adder_full fa649(.sum(ws2b4n0_21), .c_out(ws2b4n1_20), .a(ws1b6n0_21), .b(ws1b6n1_21), .c_in(wand11_31));
adder_full fa650(.sum(ws2b4n0_22), .c_out(ws2b4n1_21), .a(ws1b6n0_22), .b(ws1b6n1_22), .c_in(wand10_31));
adder_full fa651(.sum(ws2b4n0_23), .c_out(ws2b4n1_22), .a(ws1b6n0_23), .b(ws1b6n1_23), .c_in(wand9_31));
adder_full fa652(.sum(ws2b4n0_24), .c_out(ws2b4n1_23), .a(ws1b6n0_24), .b(ws1b6n1_24), .c_in(wand8_31));
adder_full fa653(.sum(ws2b4n0_25), .c_out(ws2b4n1_24), .a(ws1b6n0_25), .b(ws1b6n1_25), .c_in(wand7_31));
adder_full fa654(.sum(ws2b4n0_26), .c_out(ws2b4n1_25), .a(ws1b6n0_26), .b(ws1b6n1_26), .c_in(wand6_31));
adder_full fa655(.sum(ws2b4n0_27), .c_out(ws2b4n1_26), .a(ws1b6n0_27), .b(ws1b6n1_27), .c_in(wand5_31));
adder_full fa656(.sum(ws2b4n0_28), .c_out(ws2b4n1_27), .a(ws1b6n0_28), .b(ws1b6n1_28), .c_in(wand4_31));
adder_full fa657(.sum(ws2b4n0_29), .c_out(ws2b4n1_28), .a(ws1b6n0_29), .b(ws1b6n1_29), .c_in(wand3_31));
adder_full fa658(.sum(ws2b4n0_30), .c_out(ws2b4n1_29), .a(ws1b6n0_30), .b(ws1b6n1_30), .c_in(wand2_31));
adder_full fa659(.sum(ws2b4n0_31), .c_out(ws2b4n1_30), .a(ws1b6n0_31), .b(ws1b6n1_31), .c_in(wand1_31));
adder_full fa660(.sum(ws2b4n0_32), .c_out(ws2b4n1_31), .a(ws1b6n0_32), .b(ws1b6n1_32), .c_in(wand0_31));
adder_half ha58(.sum(ws2b4n0_33), .c_out(ws2b4n1_32), .a(ws1b6n0_33), .b(ws1b6n1_33));
assign ws2b4n0_34 = ws1b6n0_34;
assign ws2b4n0_35 = ws1b6n0_35;
assign ws2b4n0_36 = ws1b6n0_36;

assign ws3b0n0_18 = ws2b1n0_18;
assign ws3b0n0_19 = ws2b1n0_19;
assign ws3b0n0_20 = ws2b1n0_20;
assign ws3b0n0_21 = ws2b1n0_21;
assign ws3b0n0_22 = ws2b1n0_22;
assign ws3b0n0_23 = ws2b1n0_23;
adder_half ha59(.sum(ws3b0n0_24), .c_out(ws3b0n1_23), .a(ws2b0n0_24), .b(ws2b1n0_24));
adder_half ha60(.sum(ws3b0n0_25), .c_out(ws3b0n1_24), .a(ws2b0n0_25), .b(ws2b1n0_25));
adder_full fa661(.sum(ws3b0n0_26), .c_out(ws3b0n1_25), .a(ws2b0n0_26), .b(ws2b0n1_26), .c_in(ws2b1n0_26));
adder_full fa662(.sum(ws3b0n0_27), .c_out(ws3b0n1_26), .a(ws2b0n0_27), .b(ws2b0n1_27), .c_in(ws2b1n0_27));
adder_full fa663(.sum(ws3b0n0_28), .c_out(ws3b0n1_27), .a(ws2b0n0_28), .b(ws2b0n1_28), .c_in(ws2b1n0_28));
adder_full fa664(.sum(ws3b0n0_29), .c_out(ws3b0n1_28), .a(ws2b0n0_29), .b(ws2b0n1_29), .c_in(ws2b1n0_29));
adder_full fa665(.sum(ws3b0n0_30), .c_out(ws3b0n1_29), .a(ws2b0n0_30), .b(ws2b0n1_30), .c_in(ws2b1n0_30));
adder_full fa666(.sum(ws3b0n0_31), .c_out(ws3b0n1_30), .a(ws2b0n0_31), .b(ws2b0n1_31), .c_in(ws2b1n0_31));
adder_full fa667(.sum(ws3b0n0_32), .c_out(ws3b0n1_31), .a(ws2b0n0_32), .b(ws2b0n1_32), .c_in(ws2b1n0_32));
adder_full fa668(.sum(ws3b0n0_33), .c_out(ws3b0n1_32), .a(ws2b0n0_33), .b(ws2b0n1_33), .c_in(ws2b1n0_33));
adder_full fa669(.sum(ws3b0n0_34), .c_out(ws3b0n1_33), .a(ws2b0n0_34), .b(ws2b0n1_34), .c_in(ws2b1n0_34));
adder_full fa670(.sum(ws3b0n0_35), .c_out(ws3b0n1_34), .a(ws2b0n0_35), .b(ws2b0n1_35), .c_in(ws2b1n0_35));
adder_full fa671(.sum(ws3b0n0_36), .c_out(ws3b0n1_35), .a(ws2b0n0_36), .b(ws2b0n1_36), .c_in(ws2b1n0_36));
adder_full fa672(.sum(ws3b0n0_37), .c_out(ws3b0n1_36), .a(ws2b0n0_37), .b(ws2b0n1_37), .c_in(ws2b1n0_37));
adder_full fa673(.sum(ws3b0n0_38), .c_out(ws3b0n1_37), .a(ws2b0n0_38), .b(ws2b0n1_38), .c_in(ws2b1n0_38));
adder_full fa674(.sum(ws3b0n0_39), .c_out(ws3b0n1_38), .a(ws2b0n0_39), .b(ws2b0n1_39), .c_in(ws2b1n0_39));
adder_full fa675(.sum(ws3b0n0_40), .c_out(ws3b0n1_39), .a(ws2b0n0_40), .b(ws2b0n1_40), .c_in(ws2b1n0_40));
adder_full fa676(.sum(ws3b0n0_41), .c_out(ws3b0n1_40), .a(ws2b0n0_41), .b(ws2b0n1_41), .c_in(ws2b1n0_41));
adder_full fa677(.sum(ws3b0n0_42), .c_out(ws3b0n1_41), .a(ws2b0n0_42), .b(ws2b0n1_42), .c_in(ws2b1n0_42));
adder_full fa678(.sum(ws3b0n0_43), .c_out(ws3b0n1_42), .a(ws2b0n0_43), .b(ws2b0n1_43), .c_in(ws2b1n0_43));
adder_full fa679(.sum(ws3b0n0_44), .c_out(ws3b0n1_43), .a(ws2b0n0_44), .b(ws2b0n1_44), .c_in(ws2b1n0_44));
adder_full fa680(.sum(ws3b0n0_45), .c_out(ws3b0n1_44), .a(ws2b0n0_45), .b(ws2b0n1_45), .c_in(ws2b1n0_45));
adder_full fa681(.sum(ws3b0n0_46), .c_out(ws3b0n1_45), .a(ws2b0n0_46), .b(ws2b0n1_46), .c_in(ws2b1n0_46));
adder_full fa682(.sum(ws3b0n0_47), .c_out(ws3b0n1_46), .a(ws2b0n0_47), .b(ws2b0n1_47), .c_in(ws2b1n0_47));
adder_full fa683(.sum(ws3b0n0_48), .c_out(ws3b0n1_47), .a(ws2b0n0_48), .b(ws2b0n1_48), .c_in(ws2b1n0_48));
adder_full fa684(.sum(ws3b0n0_49), .c_out(ws3b0n1_48), .a(ws2b0n0_49), .b(ws2b0n1_49), .c_in(ws2b1n0_49));
adder_full fa685(.sum(ws3b0n0_50), .c_out(ws3b0n1_49), .a(ws2b0n0_50), .b(ws2b0n1_50), .c_in(ws2b1n0_50));
adder_full fa686(.sum(ws3b0n0_51), .c_out(ws3b0n1_50), .a(ws2b0n0_51), .b(ws2b0n1_51), .c_in(ws2b1n0_51));
adder_full fa687(.sum(ws3b0n0_52), .c_out(ws3b0n1_51), .a(ws2b0n0_52), .b(ws2b0n1_52), .c_in(ws2b1n0_52));
adder_full fa688(.sum(ws3b0n0_53), .c_out(ws3b0n1_52), .a(ws2b0n0_53), .b(ws2b0n1_53), .c_in(ws2b1n0_53));
adder_full fa689(.sum(ws3b0n0_54), .c_out(ws3b0n1_53), .a(ws2b0n0_54), .b(ws2b0n1_54), .c_in(ws2b1n0_54));
adder_full fa690(.sum(ws3b0n0_55), .c_out(ws3b0n1_54), .a(ws2b0n0_55), .b(ws2b0n1_55), .c_in(ws2b1n0_55));
adder_full fa691(.sum(ws3b0n0_56), .c_out(ws3b0n1_55), .a(ws2b0n0_56), .b(ws2b0n1_56), .c_in(ws2b1n0_56));
adder_half ha61(.sum(ws3b0n0_57), .c_out(ws3b0n1_56), .a(ws2b0n0_57), .b(ws2b0n1_57));
adder_half ha62(.sum(ws3b0n0_58), .c_out(ws3b0n1_57), .a(ws2b0n0_58), .b(ws2b0n1_58));
adder_half ha63(.sum(ws3b0n0_59), .c_out(ws3b0n1_58), .a(ws2b0n0_59), .b(ws2b0n1_59));
assign ws3b0n0_60 = ws2b0n0_60;
assign ws3b0n0_61 = ws2b0n0_61;
assign ws3b0n0_62 = ws2b0n0_62;
assign ws3b0n0_63 = ws2b0n0_63;
assign ws3b1n0_9 = ws2b2n0_9;
assign ws3b1n0_10 = ws2b2n0_10;
assign ws3b1n0_11 = ws2b2n0_11;
assign ws3b1n0_12 = ws2b2n0_12;
adder_half ha64(.sum(ws3b1n0_13), .c_out(ws3b1n1_12), .a(ws2b2n0_13), .b(ws2b2n1_13));
adder_half ha65(.sum(ws3b1n0_14), .c_out(ws3b1n1_13), .a(ws2b2n0_14), .b(ws2b2n1_14));
adder_half ha66(.sum(ws3b1n0_15), .c_out(ws3b1n1_14), .a(ws2b2n0_15), .b(ws2b2n1_15));
adder_half ha67(.sum(ws3b1n0_16), .c_out(ws3b1n1_15), .a(ws2b2n0_16), .b(ws2b2n1_16));
adder_half ha68(.sum(ws3b1n0_17), .c_out(ws3b1n1_16), .a(ws2b2n0_17), .b(ws2b2n1_17));
adder_half ha69(.sum(ws3b1n0_18), .c_out(ws3b1n1_17), .a(ws2b2n0_18), .b(ws2b2n1_18));
adder_full fa692(.sum(ws3b1n0_19), .c_out(ws3b1n1_18), .a(ws2b1n1_19), .b(ws2b2n0_19), .c_in(ws2b2n1_19));
adder_full fa693(.sum(ws3b1n0_20), .c_out(ws3b1n1_19), .a(ws2b1n1_20), .b(ws2b2n0_20), .c_in(ws2b2n1_20));
adder_full fa694(.sum(ws3b1n0_21), .c_out(ws3b1n1_20), .a(ws2b1n1_21), .b(ws2b2n0_21), .c_in(ws2b2n1_21));
adder_full fa695(.sum(ws3b1n0_22), .c_out(ws3b1n1_21), .a(ws2b1n1_22), .b(ws2b2n0_22), .c_in(ws2b2n1_22));
adder_full fa696(.sum(ws3b1n0_23), .c_out(ws3b1n1_22), .a(ws2b1n1_23), .b(ws2b2n0_23), .c_in(ws2b2n1_23));
adder_full fa697(.sum(ws3b1n0_24), .c_out(ws3b1n1_23), .a(ws2b1n1_24), .b(ws2b2n0_24), .c_in(ws2b2n1_24));
adder_full fa698(.sum(ws3b1n0_25), .c_out(ws3b1n1_24), .a(ws2b1n1_25), .b(ws2b2n0_25), .c_in(ws2b2n1_25));
adder_full fa699(.sum(ws3b1n0_26), .c_out(ws3b1n1_25), .a(ws2b1n1_26), .b(ws2b2n0_26), .c_in(ws2b2n1_26));
adder_full fa700(.sum(ws3b1n0_27), .c_out(ws3b1n1_26), .a(ws2b1n1_27), .b(ws2b2n0_27), .c_in(ws2b2n1_27));
adder_full fa701(.sum(ws3b1n0_28), .c_out(ws3b1n1_27), .a(ws2b1n1_28), .b(ws2b2n0_28), .c_in(ws2b2n1_28));
adder_full fa702(.sum(ws3b1n0_29), .c_out(ws3b1n1_28), .a(ws2b1n1_29), .b(ws2b2n0_29), .c_in(ws2b2n1_29));
adder_full fa703(.sum(ws3b1n0_30), .c_out(ws3b1n1_29), .a(ws2b1n1_30), .b(ws2b2n0_30), .c_in(ws2b2n1_30));
adder_full fa704(.sum(ws3b1n0_31), .c_out(ws3b1n1_30), .a(ws2b1n1_31), .b(ws2b2n0_31), .c_in(ws2b2n1_31));
adder_full fa705(.sum(ws3b1n0_32), .c_out(ws3b1n1_31), .a(ws2b1n1_32), .b(ws2b2n0_32), .c_in(ws2b2n1_32));
adder_full fa706(.sum(ws3b1n0_33), .c_out(ws3b1n1_32), .a(ws2b1n1_33), .b(ws2b2n0_33), .c_in(ws2b2n1_33));
adder_full fa707(.sum(ws3b1n0_34), .c_out(ws3b1n1_33), .a(ws2b1n1_34), .b(ws2b2n0_34), .c_in(ws2b2n1_34));
adder_full fa708(.sum(ws3b1n0_35), .c_out(ws3b1n1_34), .a(ws2b1n1_35), .b(ws2b2n0_35), .c_in(ws2b2n1_35));
adder_full fa709(.sum(ws3b1n0_36), .c_out(ws3b1n1_35), .a(ws2b1n1_36), .b(ws2b2n0_36), .c_in(ws2b2n1_36));
adder_full fa710(.sum(ws3b1n0_37), .c_out(ws3b1n1_36), .a(ws2b1n1_37), .b(ws2b2n0_37), .c_in(ws2b2n1_37));
adder_full fa711(.sum(ws3b1n0_38), .c_out(ws3b1n1_37), .a(ws2b1n1_38), .b(ws2b2n0_38), .c_in(ws2b2n1_38));
adder_full fa712(.sum(ws3b1n0_39), .c_out(ws3b1n1_38), .a(ws2b1n1_39), .b(ws2b2n0_39), .c_in(ws2b2n1_39));
adder_full fa713(.sum(ws3b1n0_40), .c_out(ws3b1n1_39), .a(ws2b1n1_40), .b(ws2b2n0_40), .c_in(ws2b2n1_40));
adder_full fa714(.sum(ws3b1n0_41), .c_out(ws3b1n1_40), .a(ws2b1n1_41), .b(ws2b2n0_41), .c_in(ws2b2n1_41));
adder_full fa715(.sum(ws3b1n0_42), .c_out(ws3b1n1_41), .a(ws2b1n1_42), .b(ws2b2n0_42), .c_in(ws2b2n1_42));
adder_full fa716(.sum(ws3b1n0_43), .c_out(ws3b1n1_42), .a(ws2b1n1_43), .b(ws2b2n0_43), .c_in(ws2b2n1_43));
adder_full fa717(.sum(ws3b1n0_44), .c_out(ws3b1n1_43), .a(ws2b1n1_44), .b(ws2b2n0_44), .c_in(ws2b2n1_44));
adder_full fa718(.sum(ws3b1n0_45), .c_out(ws3b1n1_44), .a(ws2b1n1_45), .b(ws2b2n0_45), .c_in(ws2b2n1_45));
adder_full fa719(.sum(ws3b1n0_46), .c_out(ws3b1n1_45), .a(ws2b1n1_46), .b(ws2b2n0_46), .c_in(ws2b2n1_46));
adder_half ha70(.sum(ws3b1n0_47), .c_out(ws3b1n1_46), .a(ws2b1n1_47), .b(ws2b2n0_47));
adder_half ha71(.sum(ws3b1n0_48), .c_out(ws3b1n1_47), .a(ws2b1n1_48), .b(ws2b2n0_48));
adder_half ha72(.sum(ws3b1n0_49), .c_out(ws3b1n1_48), .a(ws2b1n1_49), .b(ws2b2n0_49));
assign ws3b1n0_50 = ws2b1n1_50;
assign ws3b1n0_51 = ws2b1n1_51;
assign ws3b1n0_52 = ws2b1n1_52;
assign ws3b1n0_53 = ws2b1n1_53;
assign ws3b2n0_1 = ws2b4n0_1;
assign ws3b2n0_2 = ws2b4n0_2;
assign ws3b2n0_3 = ws2b4n0_3;
assign ws3b2n0_4 = ws2b4n0_4;
adder_full fa720(.sum(ws3b2n0_5), .c_out(ws3b2n1_4), .a(ws2b3n0_5), .b(ws2b3n1_5), .c_in(ws2b4n0_5));
adder_full fa721(.sum(ws3b2n0_6), .c_out(ws3b2n1_5), .a(ws2b3n0_6), .b(ws2b3n1_6), .c_in(ws2b4n0_6));
adder_full fa722(.sum(ws3b2n0_7), .c_out(ws3b2n1_6), .a(ws2b3n0_7), .b(ws2b3n1_7), .c_in(ws2b4n0_7));
adder_full fa723(.sum(ws3b2n0_8), .c_out(ws3b2n1_7), .a(ws2b3n0_8), .b(ws2b3n1_8), .c_in(ws2b4n0_8));
adder_full fa724(.sum(ws3b2n0_9), .c_out(ws3b2n1_8), .a(ws2b3n0_9), .b(ws2b3n1_9), .c_in(ws2b4n0_9));
adder_full fa725(.sum(ws3b2n0_10), .c_out(ws3b2n1_9), .a(ws2b3n0_10), .b(ws2b3n1_10), .c_in(ws2b4n0_10));
adder_full fa726(.sum(ws3b2n0_11), .c_out(ws3b2n1_10), .a(ws2b3n0_11), .b(ws2b3n1_11), .c_in(ws2b4n0_11));
adder_full fa727(.sum(ws3b2n0_12), .c_out(ws3b2n1_11), .a(ws2b3n0_12), .b(ws2b3n1_12), .c_in(ws2b4n0_12));
adder_full fa728(.sum(ws3b2n0_13), .c_out(ws3b2n1_12), .a(ws2b3n0_13), .b(ws2b3n1_13), .c_in(ws2b4n0_13));
adder_full fa729(.sum(ws3b2n0_14), .c_out(ws3b2n1_13), .a(ws2b3n0_14), .b(ws2b3n1_14), .c_in(ws2b4n0_14));
adder_full fa730(.sum(ws3b2n0_15), .c_out(ws3b2n1_14), .a(ws2b3n0_15), .b(ws2b3n1_15), .c_in(ws2b4n0_15));
adder_full fa731(.sum(ws3b2n0_16), .c_out(ws3b2n1_15), .a(ws2b3n0_16), .b(ws2b3n1_16), .c_in(ws2b4n0_16));
adder_full fa732(.sum(ws3b2n0_17), .c_out(ws3b2n1_16), .a(ws2b3n0_17), .b(ws2b3n1_17), .c_in(ws2b4n0_17));
adder_full fa733(.sum(ws3b2n0_18), .c_out(ws3b2n1_17), .a(ws2b3n0_18), .b(ws2b3n1_18), .c_in(ws2b4n0_18));
adder_full fa734(.sum(ws3b2n0_19), .c_out(ws3b2n1_18), .a(ws2b3n0_19), .b(ws2b3n1_19), .c_in(ws2b4n0_19));
adder_full fa735(.sum(ws3b2n0_20), .c_out(ws3b2n1_19), .a(ws2b3n0_20), .b(ws2b3n1_20), .c_in(ws2b4n0_20));
adder_full fa736(.sum(ws3b2n0_21), .c_out(ws3b2n1_20), .a(ws2b3n0_21), .b(ws2b3n1_21), .c_in(ws2b4n0_21));
adder_full fa737(.sum(ws3b2n0_22), .c_out(ws3b2n1_21), .a(ws2b3n0_22), .b(ws2b3n1_22), .c_in(ws2b4n0_22));
adder_full fa738(.sum(ws3b2n0_23), .c_out(ws3b2n1_22), .a(ws2b3n0_23), .b(ws2b3n1_23), .c_in(ws2b4n0_23));
adder_full fa739(.sum(ws3b2n0_24), .c_out(ws3b2n1_23), .a(ws2b3n0_24), .b(ws2b3n1_24), .c_in(ws2b4n0_24));
adder_full fa740(.sum(ws3b2n0_25), .c_out(ws3b2n1_24), .a(ws2b3n0_25), .b(ws2b3n1_25), .c_in(ws2b4n0_25));
adder_full fa741(.sum(ws3b2n0_26), .c_out(ws3b2n1_25), .a(ws2b3n0_26), .b(ws2b3n1_26), .c_in(ws2b4n0_26));
adder_full fa742(.sum(ws3b2n0_27), .c_out(ws3b2n1_26), .a(ws2b3n0_27), .b(ws2b3n1_27), .c_in(ws2b4n0_27));
adder_full fa743(.sum(ws3b2n0_28), .c_out(ws3b2n1_27), .a(ws2b3n0_28), .b(ws2b3n1_28), .c_in(ws2b4n0_28));
adder_full fa744(.sum(ws3b2n0_29), .c_out(ws3b2n1_28), .a(ws2b3n0_29), .b(ws2b3n1_29), .c_in(ws2b4n0_29));
adder_full fa745(.sum(ws3b2n0_30), .c_out(ws3b2n1_29), .a(ws2b3n0_30), .b(ws2b3n1_30), .c_in(ws2b4n0_30));
adder_full fa746(.sum(ws3b2n0_31), .c_out(ws3b2n1_30), .a(ws2b3n0_31), .b(ws2b3n1_31), .c_in(ws2b4n0_31));
adder_full fa747(.sum(ws3b2n0_32), .c_out(ws3b2n1_31), .a(ws2b3n0_32), .b(ws2b3n1_32), .c_in(ws2b4n0_32));
adder_full fa748(.sum(ws3b2n0_33), .c_out(ws3b2n1_32), .a(ws2b3n0_33), .b(ws2b3n1_33), .c_in(ws2b4n0_33));
adder_full fa749(.sum(ws3b2n0_34), .c_out(ws3b2n1_33), .a(ws2b3n0_34), .b(ws2b3n1_34), .c_in(ws2b4n0_34));
adder_full fa750(.sum(ws3b2n0_35), .c_out(ws3b2n1_34), .a(ws2b3n0_35), .b(ws2b3n1_35), .c_in(ws2b4n0_35));
adder_full fa751(.sum(ws3b2n0_36), .c_out(ws3b2n1_35), .a(ws2b3n0_36), .b(ws2b3n1_36), .c_in(ws2b4n0_36));
adder_half ha73(.sum(ws3b2n0_37), .c_out(ws3b2n1_36), .a(ws2b3n0_37), .b(ws2b3n1_37));
adder_half ha74(.sum(ws3b2n0_38), .c_out(ws3b2n1_37), .a(ws2b3n0_38), .b(ws2b3n1_38));
adder_half ha75(.sum(ws3b2n0_39), .c_out(ws3b2n1_38), .a(ws2b3n0_39), .b(ws2b3n1_39));
assign ws3b2n0_40 = ws2b3n0_40;
assign ws3b2n0_41 = ws2b3n0_41;
assign ws3b2n0_42 = ws2b3n0_42;

assign ws4b0n0_9 = ws3b1n0_9;
assign ws4b0n0_10 = ws3b1n0_10;
assign ws4b0n0_11 = ws3b1n0_11;
assign ws4b0n0_12 = ws3b1n0_12;
assign ws4b0n0_13 = ws3b1n0_13;
assign ws4b0n0_14 = ws3b1n0_14;
assign ws4b0n0_15 = ws3b1n0_15;
assign ws4b0n0_16 = ws3b1n0_16;
assign ws4b0n0_17 = ws3b1n0_17;
adder_half ha76(.sum(ws4b0n0_18), .c_out(ws4b0n1_17), .a(ws3b0n0_18), .b(ws3b1n0_18));
adder_half ha77(.sum(ws4b0n0_19), .c_out(ws4b0n1_18), .a(ws3b0n0_19), .b(ws3b1n0_19));
adder_half ha78(.sum(ws4b0n0_20), .c_out(ws4b0n1_19), .a(ws3b0n0_20), .b(ws3b1n0_20));
adder_half ha79(.sum(ws4b0n0_21), .c_out(ws4b0n1_20), .a(ws3b0n0_21), .b(ws3b1n0_21));
adder_half ha80(.sum(ws4b0n0_22), .c_out(ws4b0n1_21), .a(ws3b0n0_22), .b(ws3b1n0_22));
adder_full fa752(.sum(ws4b0n0_23), .c_out(ws4b0n1_22), .a(ws3b0n0_23), .b(ws3b0n1_23), .c_in(ws3b1n0_23));
adder_full fa753(.sum(ws4b0n0_24), .c_out(ws4b0n1_23), .a(ws3b0n0_24), .b(ws3b0n1_24), .c_in(ws3b1n0_24));
adder_full fa754(.sum(ws4b0n0_25), .c_out(ws4b0n1_24), .a(ws3b0n0_25), .b(ws3b0n1_25), .c_in(ws3b1n0_25));
adder_full fa755(.sum(ws4b0n0_26), .c_out(ws4b0n1_25), .a(ws3b0n0_26), .b(ws3b0n1_26), .c_in(ws3b1n0_26));
adder_full fa756(.sum(ws4b0n0_27), .c_out(ws4b0n1_26), .a(ws3b0n0_27), .b(ws3b0n1_27), .c_in(ws3b1n0_27));
adder_full fa757(.sum(ws4b0n0_28), .c_out(ws4b0n1_27), .a(ws3b0n0_28), .b(ws3b0n1_28), .c_in(ws3b1n0_28));
adder_full fa758(.sum(ws4b0n0_29), .c_out(ws4b0n1_28), .a(ws3b0n0_29), .b(ws3b0n1_29), .c_in(ws3b1n0_29));
adder_full fa759(.sum(ws4b0n0_30), .c_out(ws4b0n1_29), .a(ws3b0n0_30), .b(ws3b0n1_30), .c_in(ws3b1n0_30));
adder_full fa760(.sum(ws4b0n0_31), .c_out(ws4b0n1_30), .a(ws3b0n0_31), .b(ws3b0n1_31), .c_in(ws3b1n0_31));
adder_full fa761(.sum(ws4b0n0_32), .c_out(ws4b0n1_31), .a(ws3b0n0_32), .b(ws3b0n1_32), .c_in(ws3b1n0_32));
adder_full fa762(.sum(ws4b0n0_33), .c_out(ws4b0n1_32), .a(ws3b0n0_33), .b(ws3b0n1_33), .c_in(ws3b1n0_33));
adder_full fa763(.sum(ws4b0n0_34), .c_out(ws4b0n1_33), .a(ws3b0n0_34), .b(ws3b0n1_34), .c_in(ws3b1n0_34));
adder_full fa764(.sum(ws4b0n0_35), .c_out(ws4b0n1_34), .a(ws3b0n0_35), .b(ws3b0n1_35), .c_in(ws3b1n0_35));
adder_full fa765(.sum(ws4b0n0_36), .c_out(ws4b0n1_35), .a(ws3b0n0_36), .b(ws3b0n1_36), .c_in(ws3b1n0_36));
adder_full fa766(.sum(ws4b0n0_37), .c_out(ws4b0n1_36), .a(ws3b0n0_37), .b(ws3b0n1_37), .c_in(ws3b1n0_37));
adder_full fa767(.sum(ws4b0n0_38), .c_out(ws4b0n1_37), .a(ws3b0n0_38), .b(ws3b0n1_38), .c_in(ws3b1n0_38));
adder_full fa768(.sum(ws4b0n0_39), .c_out(ws4b0n1_38), .a(ws3b0n0_39), .b(ws3b0n1_39), .c_in(ws3b1n0_39));
adder_full fa769(.sum(ws4b0n0_40), .c_out(ws4b0n1_39), .a(ws3b0n0_40), .b(ws3b0n1_40), .c_in(ws3b1n0_40));
adder_full fa770(.sum(ws4b0n0_41), .c_out(ws4b0n1_40), .a(ws3b0n0_41), .b(ws3b0n1_41), .c_in(ws3b1n0_41));
adder_full fa771(.sum(ws4b0n0_42), .c_out(ws4b0n1_41), .a(ws3b0n0_42), .b(ws3b0n1_42), .c_in(ws3b1n0_42));
adder_full fa772(.sum(ws4b0n0_43), .c_out(ws4b0n1_42), .a(ws3b0n0_43), .b(ws3b0n1_43), .c_in(ws3b1n0_43));
adder_full fa773(.sum(ws4b0n0_44), .c_out(ws4b0n1_43), .a(ws3b0n0_44), .b(ws3b0n1_44), .c_in(ws3b1n0_44));
adder_full fa774(.sum(ws4b0n0_45), .c_out(ws4b0n1_44), .a(ws3b0n0_45), .b(ws3b0n1_45), .c_in(ws3b1n0_45));
adder_full fa775(.sum(ws4b0n0_46), .c_out(ws4b0n1_45), .a(ws3b0n0_46), .b(ws3b0n1_46), .c_in(ws3b1n0_46));
adder_full fa776(.sum(ws4b0n0_47), .c_out(ws4b0n1_46), .a(ws3b0n0_47), .b(ws3b0n1_47), .c_in(ws3b1n0_47));
adder_full fa777(.sum(ws4b0n0_48), .c_out(ws4b0n1_47), .a(ws3b0n0_48), .b(ws3b0n1_48), .c_in(ws3b1n0_48));
adder_full fa778(.sum(ws4b0n0_49), .c_out(ws4b0n1_48), .a(ws3b0n0_49), .b(ws3b0n1_49), .c_in(ws3b1n0_49));
adder_full fa779(.sum(ws4b0n0_50), .c_out(ws4b0n1_49), .a(ws3b0n0_50), .b(ws3b0n1_50), .c_in(ws3b1n0_50));
adder_full fa780(.sum(ws4b0n0_51), .c_out(ws4b0n1_50), .a(ws3b0n0_51), .b(ws3b0n1_51), .c_in(ws3b1n0_51));
adder_full fa781(.sum(ws4b0n0_52), .c_out(ws4b0n1_51), .a(ws3b0n0_52), .b(ws3b0n1_52), .c_in(ws3b1n0_52));
adder_full fa782(.sum(ws4b0n0_53), .c_out(ws4b0n1_52), .a(ws3b0n0_53), .b(ws3b0n1_53), .c_in(ws3b1n0_53));
adder_half ha81(.sum(ws4b0n0_54), .c_out(ws4b0n1_53), .a(ws3b0n0_54), .b(ws3b0n1_54));
adder_half ha82(.sum(ws4b0n0_55), .c_out(ws4b0n1_54), .a(ws3b0n0_55), .b(ws3b0n1_55));
adder_half ha83(.sum(ws4b0n0_56), .c_out(ws4b0n1_55), .a(ws3b0n0_56), .b(ws3b0n1_56));
adder_half ha84(.sum(ws4b0n0_57), .c_out(ws4b0n1_56), .a(ws3b0n0_57), .b(ws3b0n1_57));
adder_half ha85(.sum(ws4b0n0_58), .c_out(ws4b0n1_57), .a(ws3b0n0_58), .b(ws3b0n1_58));
assign ws4b0n0_59 = ws3b0n0_59;
assign ws4b0n0_60 = ws3b0n0_60;
assign ws4b0n0_61 = ws3b0n0_61;
assign ws4b0n0_62 = ws3b0n0_62;
assign ws4b0n0_63 = ws3b0n0_63;
assign ws4b1n0_1 = ws3b2n0_1;
assign ws4b1n0_2 = ws3b2n0_2;
assign ws4b1n0_3 = ws3b2n0_3;
adder_half ha86(.sum(ws4b1n0_4), .c_out(ws4b1n1_3), .a(ws3b2n0_4), .b(ws3b2n1_4));
adder_half ha87(.sum(ws4b1n0_5), .c_out(ws4b1n1_4), .a(ws3b2n0_5), .b(ws3b2n1_5));
adder_half ha88(.sum(ws4b1n0_6), .c_out(ws4b1n1_5), .a(ws3b2n0_6), .b(ws3b2n1_6));
adder_half ha89(.sum(ws4b1n0_7), .c_out(ws4b1n1_6), .a(ws3b2n0_7), .b(ws3b2n1_7));
adder_half ha90(.sum(ws4b1n0_8), .c_out(ws4b1n1_7), .a(ws3b2n0_8), .b(ws3b2n1_8));
adder_half ha91(.sum(ws4b1n0_9), .c_out(ws4b1n1_8), .a(ws3b2n0_9), .b(ws3b2n1_9));
adder_half ha92(.sum(ws4b1n0_10), .c_out(ws4b1n1_9), .a(ws3b2n0_10), .b(ws3b2n1_10));
adder_half ha93(.sum(ws4b1n0_11), .c_out(ws4b1n1_10), .a(ws3b2n0_11), .b(ws3b2n1_11));
adder_full fa783(.sum(ws4b1n0_12), .c_out(ws4b1n1_11), .a(ws3b1n1_12), .b(ws3b2n0_12), .c_in(ws3b2n1_12));
adder_full fa784(.sum(ws4b1n0_13), .c_out(ws4b1n1_12), .a(ws3b1n1_13), .b(ws3b2n0_13), .c_in(ws3b2n1_13));
adder_full fa785(.sum(ws4b1n0_14), .c_out(ws4b1n1_13), .a(ws3b1n1_14), .b(ws3b2n0_14), .c_in(ws3b2n1_14));
adder_full fa786(.sum(ws4b1n0_15), .c_out(ws4b1n1_14), .a(ws3b1n1_15), .b(ws3b2n0_15), .c_in(ws3b2n1_15));
adder_full fa787(.sum(ws4b1n0_16), .c_out(ws4b1n1_15), .a(ws3b1n1_16), .b(ws3b2n0_16), .c_in(ws3b2n1_16));
adder_full fa788(.sum(ws4b1n0_17), .c_out(ws4b1n1_16), .a(ws3b1n1_17), .b(ws3b2n0_17), .c_in(ws3b2n1_17));
adder_full fa789(.sum(ws4b1n0_18), .c_out(ws4b1n1_17), .a(ws3b1n1_18), .b(ws3b2n0_18), .c_in(ws3b2n1_18));
adder_full fa790(.sum(ws4b1n0_19), .c_out(ws4b1n1_18), .a(ws3b1n1_19), .b(ws3b2n0_19), .c_in(ws3b2n1_19));
adder_full fa791(.sum(ws4b1n0_20), .c_out(ws4b1n1_19), .a(ws3b1n1_20), .b(ws3b2n0_20), .c_in(ws3b2n1_20));
adder_full fa792(.sum(ws4b1n0_21), .c_out(ws4b1n1_20), .a(ws3b1n1_21), .b(ws3b2n0_21), .c_in(ws3b2n1_21));
adder_full fa793(.sum(ws4b1n0_22), .c_out(ws4b1n1_21), .a(ws3b1n1_22), .b(ws3b2n0_22), .c_in(ws3b2n1_22));
adder_full fa794(.sum(ws4b1n0_23), .c_out(ws4b1n1_22), .a(ws3b1n1_23), .b(ws3b2n0_23), .c_in(ws3b2n1_23));
adder_full fa795(.sum(ws4b1n0_24), .c_out(ws4b1n1_23), .a(ws3b1n1_24), .b(ws3b2n0_24), .c_in(ws3b2n1_24));
adder_full fa796(.sum(ws4b1n0_25), .c_out(ws4b1n1_24), .a(ws3b1n1_25), .b(ws3b2n0_25), .c_in(ws3b2n1_25));
adder_full fa797(.sum(ws4b1n0_26), .c_out(ws4b1n1_25), .a(ws3b1n1_26), .b(ws3b2n0_26), .c_in(ws3b2n1_26));
adder_full fa798(.sum(ws4b1n0_27), .c_out(ws4b1n1_26), .a(ws3b1n1_27), .b(ws3b2n0_27), .c_in(ws3b2n1_27));
adder_full fa799(.sum(ws4b1n0_28), .c_out(ws4b1n1_27), .a(ws3b1n1_28), .b(ws3b2n0_28), .c_in(ws3b2n1_28));
adder_full fa800(.sum(ws4b1n0_29), .c_out(ws4b1n1_28), .a(ws3b1n1_29), .b(ws3b2n0_29), .c_in(ws3b2n1_29));
adder_full fa801(.sum(ws4b1n0_30), .c_out(ws4b1n1_29), .a(ws3b1n1_30), .b(ws3b2n0_30), .c_in(ws3b2n1_30));
adder_full fa802(.sum(ws4b1n0_31), .c_out(ws4b1n1_30), .a(ws3b1n1_31), .b(ws3b2n0_31), .c_in(ws3b2n1_31));
adder_full fa803(.sum(ws4b1n0_32), .c_out(ws4b1n1_31), .a(ws3b1n1_32), .b(ws3b2n0_32), .c_in(ws3b2n1_32));
adder_full fa804(.sum(ws4b1n0_33), .c_out(ws4b1n1_32), .a(ws3b1n1_33), .b(ws3b2n0_33), .c_in(ws3b2n1_33));
adder_full fa805(.sum(ws4b1n0_34), .c_out(ws4b1n1_33), .a(ws3b1n1_34), .b(ws3b2n0_34), .c_in(ws3b2n1_34));
adder_full fa806(.sum(ws4b1n0_35), .c_out(ws4b1n1_34), .a(ws3b1n1_35), .b(ws3b2n0_35), .c_in(ws3b2n1_35));
adder_full fa807(.sum(ws4b1n0_36), .c_out(ws4b1n1_35), .a(ws3b1n1_36), .b(ws3b2n0_36), .c_in(ws3b2n1_36));
adder_full fa808(.sum(ws4b1n0_37), .c_out(ws4b1n1_36), .a(ws3b1n1_37), .b(ws3b2n0_37), .c_in(ws3b2n1_37));
adder_full fa809(.sum(ws4b1n0_38), .c_out(ws4b1n1_37), .a(ws3b1n1_38), .b(ws3b2n0_38), .c_in(ws3b2n1_38));
adder_half ha94(.sum(ws4b1n0_39), .c_out(ws4b1n1_38), .a(ws3b1n1_39), .b(ws3b2n0_39));
adder_half ha95(.sum(ws4b1n0_40), .c_out(ws4b1n1_39), .a(ws3b1n1_40), .b(ws3b2n0_40));
adder_half ha96(.sum(ws4b1n0_41), .c_out(ws4b1n1_40), .a(ws3b1n1_41), .b(ws3b2n0_41));
adder_half ha97(.sum(ws4b1n0_42), .c_out(ws4b1n1_41), .a(ws3b1n1_42), .b(ws3b2n0_42));
assign ws4b1n0_43 = ws3b1n1_43;
assign ws4b1n0_44 = ws3b1n1_44;
assign ws4b1n0_45 = ws3b1n1_45;
assign ws4b1n0_46 = ws3b1n1_46;
assign ws4b1n0_47 = ws3b1n1_47;
assign ws4b1n0_48 = ws3b1n1_48;

assign ws5b0n0_1 = ws4b1n0_1;
assign ws5b0n0_2 = ws4b1n0_2;
assign ws5b0n0_3 = ws4b1n0_3;
assign ws5b0n0_4 = ws4b1n0_4;
assign ws5b0n0_5 = ws4b1n0_5;
assign ws5b0n0_6 = ws4b1n0_6;
assign ws5b0n0_7 = ws4b1n0_7;
assign ws5b0n0_8 = ws4b1n0_8;
adder_half ha98(.sum(ws5b0n0_9), .c_out(ws5b0n1_8), .a(ws4b0n0_9), .b(ws4b1n0_9));
adder_half ha99(.sum(ws5b0n0_10), .c_out(ws5b0n1_9), .a(ws4b0n0_10), .b(ws4b1n0_10));
adder_half ha100(.sum(ws5b0n0_11), .c_out(ws5b0n1_10), .a(ws4b0n0_11), .b(ws4b1n0_11));
adder_half ha101(.sum(ws5b0n0_12), .c_out(ws5b0n1_11), .a(ws4b0n0_12), .b(ws4b1n0_12));
adder_half ha102(.sum(ws5b0n0_13), .c_out(ws5b0n1_12), .a(ws4b0n0_13), .b(ws4b1n0_13));
adder_half ha103(.sum(ws5b0n0_14), .c_out(ws5b0n1_13), .a(ws4b0n0_14), .b(ws4b1n0_14));
adder_half ha104(.sum(ws5b0n0_15), .c_out(ws5b0n1_14), .a(ws4b0n0_15), .b(ws4b1n0_15));
adder_half ha105(.sum(ws5b0n0_16), .c_out(ws5b0n1_15), .a(ws4b0n0_16), .b(ws4b1n0_16));
adder_full fa810(.sum(ws5b0n0_17), .c_out(ws5b0n1_16), .a(ws4b0n0_17), .b(ws4b0n1_17), .c_in(ws4b1n0_17));
adder_full fa811(.sum(ws5b0n0_18), .c_out(ws5b0n1_17), .a(ws4b0n0_18), .b(ws4b0n1_18), .c_in(ws4b1n0_18));
adder_full fa812(.sum(ws5b0n0_19), .c_out(ws5b0n1_18), .a(ws4b0n0_19), .b(ws4b0n1_19), .c_in(ws4b1n0_19));
adder_full fa813(.sum(ws5b0n0_20), .c_out(ws5b0n1_19), .a(ws4b0n0_20), .b(ws4b0n1_20), .c_in(ws4b1n0_20));
adder_full fa814(.sum(ws5b0n0_21), .c_out(ws5b0n1_20), .a(ws4b0n0_21), .b(ws4b0n1_21), .c_in(ws4b1n0_21));
adder_full fa815(.sum(ws5b0n0_22), .c_out(ws5b0n1_21), .a(ws4b0n0_22), .b(ws4b0n1_22), .c_in(ws4b1n0_22));
adder_full fa816(.sum(ws5b0n0_23), .c_out(ws5b0n1_22), .a(ws4b0n0_23), .b(ws4b0n1_23), .c_in(ws4b1n0_23));
adder_full fa817(.sum(ws5b0n0_24), .c_out(ws5b0n1_23), .a(ws4b0n0_24), .b(ws4b0n1_24), .c_in(ws4b1n0_24));
adder_full fa818(.sum(ws5b0n0_25), .c_out(ws5b0n1_24), .a(ws4b0n0_25), .b(ws4b0n1_25), .c_in(ws4b1n0_25));
adder_full fa819(.sum(ws5b0n0_26), .c_out(ws5b0n1_25), .a(ws4b0n0_26), .b(ws4b0n1_26), .c_in(ws4b1n0_26));
adder_full fa820(.sum(ws5b0n0_27), .c_out(ws5b0n1_26), .a(ws4b0n0_27), .b(ws4b0n1_27), .c_in(ws4b1n0_27));
adder_full fa821(.sum(ws5b0n0_28), .c_out(ws5b0n1_27), .a(ws4b0n0_28), .b(ws4b0n1_28), .c_in(ws4b1n0_28));
adder_full fa822(.sum(ws5b0n0_29), .c_out(ws5b0n1_28), .a(ws4b0n0_29), .b(ws4b0n1_29), .c_in(ws4b1n0_29));
adder_full fa823(.sum(ws5b0n0_30), .c_out(ws5b0n1_29), .a(ws4b0n0_30), .b(ws4b0n1_30), .c_in(ws4b1n0_30));
adder_full fa824(.sum(ws5b0n0_31), .c_out(ws5b0n1_30), .a(ws4b0n0_31), .b(ws4b0n1_31), .c_in(ws4b1n0_31));
adder_full fa825(.sum(ws5b0n0_32), .c_out(ws5b0n1_31), .a(ws4b0n0_32), .b(ws4b0n1_32), .c_in(ws4b1n0_32));
adder_full fa826(.sum(ws5b0n0_33), .c_out(ws5b0n1_32), .a(ws4b0n0_33), .b(ws4b0n1_33), .c_in(ws4b1n0_33));
adder_full fa827(.sum(ws5b0n0_34), .c_out(ws5b0n1_33), .a(ws4b0n0_34), .b(ws4b0n1_34), .c_in(ws4b1n0_34));
adder_full fa828(.sum(ws5b0n0_35), .c_out(ws5b0n1_34), .a(ws4b0n0_35), .b(ws4b0n1_35), .c_in(ws4b1n0_35));
adder_full fa829(.sum(ws5b0n0_36), .c_out(ws5b0n1_35), .a(ws4b0n0_36), .b(ws4b0n1_36), .c_in(ws4b1n0_36));
adder_full fa830(.sum(ws5b0n0_37), .c_out(ws5b0n1_36), .a(ws4b0n0_37), .b(ws4b0n1_37), .c_in(ws4b1n0_37));
adder_full fa831(.sum(ws5b0n0_38), .c_out(ws5b0n1_37), .a(ws4b0n0_38), .b(ws4b0n1_38), .c_in(ws4b1n0_38));
adder_full fa832(.sum(ws5b0n0_39), .c_out(ws5b0n1_38), .a(ws4b0n0_39), .b(ws4b0n1_39), .c_in(ws4b1n0_39));
adder_full fa833(.sum(ws5b0n0_40), .c_out(ws5b0n1_39), .a(ws4b0n0_40), .b(ws4b0n1_40), .c_in(ws4b1n0_40));
adder_full fa834(.sum(ws5b0n0_41), .c_out(ws5b0n1_40), .a(ws4b0n0_41), .b(ws4b0n1_41), .c_in(ws4b1n0_41));
adder_full fa835(.sum(ws5b0n0_42), .c_out(ws5b0n1_41), .a(ws4b0n0_42), .b(ws4b0n1_42), .c_in(ws4b1n0_42));
adder_full fa836(.sum(ws5b0n0_43), .c_out(ws5b0n1_42), .a(ws4b0n0_43), .b(ws4b0n1_43), .c_in(ws4b1n0_43));
adder_full fa837(.sum(ws5b0n0_44), .c_out(ws5b0n1_43), .a(ws4b0n0_44), .b(ws4b0n1_44), .c_in(ws4b1n0_44));
adder_full fa838(.sum(ws5b0n0_45), .c_out(ws5b0n1_44), .a(ws4b0n0_45), .b(ws4b0n1_45), .c_in(ws4b1n0_45));
adder_full fa839(.sum(ws5b0n0_46), .c_out(ws5b0n1_45), .a(ws4b0n0_46), .b(ws4b0n1_46), .c_in(ws4b1n0_46));
adder_full fa840(.sum(ws5b0n0_47), .c_out(ws5b0n1_46), .a(ws4b0n0_47), .b(ws4b0n1_47), .c_in(ws4b1n0_47));
adder_full fa841(.sum(ws5b0n0_48), .c_out(ws5b0n1_47), .a(ws4b0n0_48), .b(ws4b0n1_48), .c_in(ws4b1n0_48));
adder_half ha106(.sum(ws5b0n0_49), .c_out(ws5b0n1_48), .a(ws4b0n0_49), .b(ws4b0n1_49));
adder_half ha107(.sum(ws5b0n0_50), .c_out(ws5b0n1_49), .a(ws4b0n0_50), .b(ws4b0n1_50));
adder_half ha108(.sum(ws5b0n0_51), .c_out(ws5b0n1_50), .a(ws4b0n0_51), .b(ws4b0n1_51));
adder_half ha109(.sum(ws5b0n0_52), .c_out(ws5b0n1_51), .a(ws4b0n0_52), .b(ws4b0n1_52));
adder_half ha110(.sum(ws5b0n0_53), .c_out(ws5b0n1_52), .a(ws4b0n0_53), .b(ws4b0n1_53));
adder_half ha111(.sum(ws5b0n0_54), .c_out(ws5b0n1_53), .a(ws4b0n0_54), .b(ws4b0n1_54));
adder_half ha112(.sum(ws5b0n0_55), .c_out(ws5b0n1_54), .a(ws4b0n0_55), .b(ws4b0n1_55));
adder_half ha113(.sum(ws5b0n0_56), .c_out(ws5b0n1_55), .a(ws4b0n0_56), .b(ws4b0n1_56));
adder_half ha114(.sum(ws5b0n0_57), .c_out(ws5b0n1_56), .a(ws4b0n0_57), .b(ws4b0n1_57));
assign ws5b0n0_58 = ws4b0n0_58;
assign ws5b0n0_59 = ws4b0n0_59;
assign ws5b0n0_60 = ws4b0n0_60;
assign ws5b0n0_61 = ws4b0n0_61;
assign ws5b0n0_62 = ws4b0n0_62;
assign ws5b0n0_63 = ws4b0n0_63;

assign ws6b0n0_1 = ws5b0n0_1;
assign ws6b0n0_2 = ws5b0n0_2;
adder_half ha115(.sum(ws6b0n0_3), .c_out(ws6b0n1_2), .a(ws5b0n0_3), .b(ws4b1n1_3));
adder_half ha116(.sum(ws6b0n0_4), .c_out(ws6b0n1_3), .a(ws5b0n0_4), .b(ws4b1n1_4));
adder_half ha117(.sum(ws6b0n0_5), .c_out(ws6b0n1_4), .a(ws5b0n0_5), .b(ws4b1n1_5));
adder_half ha118(.sum(ws6b0n0_6), .c_out(ws6b0n1_5), .a(ws5b0n0_6), .b(ws4b1n1_6));
adder_half ha119(.sum(ws6b0n0_7), .c_out(ws6b0n1_6), .a(ws5b0n0_7), .b(ws4b1n1_7));
adder_full fa842(.sum(ws6b0n0_8), .c_out(ws6b0n1_7), .a(ws5b0n0_8), .b(ws5b0n1_8), .c_in(ws4b1n1_8));
adder_full fa843(.sum(ws6b0n0_9), .c_out(ws6b0n1_8), .a(ws5b0n0_9), .b(ws5b0n1_9), .c_in(ws4b1n1_9));
adder_full fa844(.sum(ws6b0n0_10), .c_out(ws6b0n1_9), .a(ws5b0n0_10), .b(ws5b0n1_10), .c_in(ws4b1n1_10));
adder_full fa845(.sum(ws6b0n0_11), .c_out(ws6b0n1_10), .a(ws5b0n0_11), .b(ws5b0n1_11), .c_in(ws4b1n1_11));
adder_full fa846(.sum(ws6b0n0_12), .c_out(ws6b0n1_11), .a(ws5b0n0_12), .b(ws5b0n1_12), .c_in(ws4b1n1_12));
adder_full fa847(.sum(ws6b0n0_13), .c_out(ws6b0n1_12), .a(ws5b0n0_13), .b(ws5b0n1_13), .c_in(ws4b1n1_13));
adder_full fa848(.sum(ws6b0n0_14), .c_out(ws6b0n1_13), .a(ws5b0n0_14), .b(ws5b0n1_14), .c_in(ws4b1n1_14));
adder_full fa849(.sum(ws6b0n0_15), .c_out(ws6b0n1_14), .a(ws5b0n0_15), .b(ws5b0n1_15), .c_in(ws4b1n1_15));
adder_full fa850(.sum(ws6b0n0_16), .c_out(ws6b0n1_15), .a(ws5b0n0_16), .b(ws5b0n1_16), .c_in(ws4b1n1_16));
adder_full fa851(.sum(ws6b0n0_17), .c_out(ws6b0n1_16), .a(ws5b0n0_17), .b(ws5b0n1_17), .c_in(ws4b1n1_17));
adder_full fa852(.sum(ws6b0n0_18), .c_out(ws6b0n1_17), .a(ws5b0n0_18), .b(ws5b0n1_18), .c_in(ws4b1n1_18));
adder_full fa853(.sum(ws6b0n0_19), .c_out(ws6b0n1_18), .a(ws5b0n0_19), .b(ws5b0n1_19), .c_in(ws4b1n1_19));
adder_full fa854(.sum(ws6b0n0_20), .c_out(ws6b0n1_19), .a(ws5b0n0_20), .b(ws5b0n1_20), .c_in(ws4b1n1_20));
adder_full fa855(.sum(ws6b0n0_21), .c_out(ws6b0n1_20), .a(ws5b0n0_21), .b(ws5b0n1_21), .c_in(ws4b1n1_21));
adder_full fa856(.sum(ws6b0n0_22), .c_out(ws6b0n1_21), .a(ws5b0n0_22), .b(ws5b0n1_22), .c_in(ws4b1n1_22));
adder_full fa857(.sum(ws6b0n0_23), .c_out(ws6b0n1_22), .a(ws5b0n0_23), .b(ws5b0n1_23), .c_in(ws4b1n1_23));
adder_full fa858(.sum(ws6b0n0_24), .c_out(ws6b0n1_23), .a(ws5b0n0_24), .b(ws5b0n1_24), .c_in(ws4b1n1_24));
adder_full fa859(.sum(ws6b0n0_25), .c_out(ws6b0n1_24), .a(ws5b0n0_25), .b(ws5b0n1_25), .c_in(ws4b1n1_25));
adder_full fa860(.sum(ws6b0n0_26), .c_out(ws6b0n1_25), .a(ws5b0n0_26), .b(ws5b0n1_26), .c_in(ws4b1n1_26));
adder_full fa861(.sum(ws6b0n0_27), .c_out(ws6b0n1_26), .a(ws5b0n0_27), .b(ws5b0n1_27), .c_in(ws4b1n1_27));
adder_full fa862(.sum(ws6b0n0_28), .c_out(ws6b0n1_27), .a(ws5b0n0_28), .b(ws5b0n1_28), .c_in(ws4b1n1_28));
adder_full fa863(.sum(ws6b0n0_29), .c_out(ws6b0n1_28), .a(ws5b0n0_29), .b(ws5b0n1_29), .c_in(ws4b1n1_29));
adder_full fa864(.sum(ws6b0n0_30), .c_out(ws6b0n1_29), .a(ws5b0n0_30), .b(ws5b0n1_30), .c_in(ws4b1n1_30));
adder_full fa865(.sum(ws6b0n0_31), .c_out(ws6b0n1_30), .a(ws5b0n0_31), .b(ws5b0n1_31), .c_in(ws4b1n1_31));
adder_full fa866(.sum(ws6b0n0_32), .c_out(ws6b0n1_31), .a(ws5b0n0_32), .b(ws5b0n1_32), .c_in(ws4b1n1_32));
adder_full fa867(.sum(ws6b0n0_33), .c_out(ws6b0n1_32), .a(ws5b0n0_33), .b(ws5b0n1_33), .c_in(ws4b1n1_33));
adder_full fa868(.sum(ws6b0n0_34), .c_out(ws6b0n1_33), .a(ws5b0n0_34), .b(ws5b0n1_34), .c_in(ws4b1n1_34));
adder_full fa869(.sum(ws6b0n0_35), .c_out(ws6b0n1_34), .a(ws5b0n0_35), .b(ws5b0n1_35), .c_in(ws4b1n1_35));
adder_full fa870(.sum(ws6b0n0_36), .c_out(ws6b0n1_35), .a(ws5b0n0_36), .b(ws5b0n1_36), .c_in(ws4b1n1_36));
adder_full fa871(.sum(ws6b0n0_37), .c_out(ws6b0n1_36), .a(ws5b0n0_37), .b(ws5b0n1_37), .c_in(ws4b1n1_37));
adder_full fa872(.sum(ws6b0n0_38), .c_out(ws6b0n1_37), .a(ws5b0n0_38), .b(ws5b0n1_38), .c_in(ws4b1n1_38));
adder_full fa873(.sum(ws6b0n0_39), .c_out(ws6b0n1_38), .a(ws5b0n0_39), .b(ws5b0n1_39), .c_in(ws4b1n1_39));
adder_full fa874(.sum(ws6b0n0_40), .c_out(ws6b0n1_39), .a(ws5b0n0_40), .b(ws5b0n1_40), .c_in(ws4b1n1_40));
adder_full fa875(.sum(ws6b0n0_41), .c_out(ws6b0n1_40), .a(ws5b0n0_41), .b(ws5b0n1_41), .c_in(ws4b1n1_41));
adder_half ha120(.sum(ws6b0n0_42), .c_out(ws6b0n1_41), .a(ws5b0n0_42), .b(ws5b0n1_42));
adder_half ha121(.sum(ws6b0n0_43), .c_out(ws6b0n1_42), .a(ws5b0n0_43), .b(ws5b0n1_43));
adder_half ha122(.sum(ws6b0n0_44), .c_out(ws6b0n1_43), .a(ws5b0n0_44), .b(ws5b0n1_44));
adder_half ha123(.sum(ws6b0n0_45), .c_out(ws6b0n1_44), .a(ws5b0n0_45), .b(ws5b0n1_45));
adder_half ha124(.sum(ws6b0n0_46), .c_out(ws6b0n1_45), .a(ws5b0n0_46), .b(ws5b0n1_46));
adder_half ha125(.sum(ws6b0n0_47), .c_out(ws6b0n1_46), .a(ws5b0n0_47), .b(ws5b0n1_47));
adder_half ha126(.sum(ws6b0n0_48), .c_out(ws6b0n1_47), .a(ws5b0n0_48), .b(ws5b0n1_48));
adder_half ha127(.sum(ws6b0n0_49), .c_out(ws6b0n1_48), .a(ws5b0n0_49), .b(ws5b0n1_49));
adder_half ha128(.sum(ws6b0n0_50), .c_out(ws6b0n1_49), .a(ws5b0n0_50), .b(ws5b0n1_50));
adder_half ha129(.sum(ws6b0n0_51), .c_out(ws6b0n1_50), .a(ws5b0n0_51), .b(ws5b0n1_51));
adder_half ha130(.sum(ws6b0n0_52), .c_out(ws6b0n1_51), .a(ws5b0n0_52), .b(ws5b0n1_52));
adder_half ha131(.sum(ws6b0n0_53), .c_out(ws6b0n1_52), .a(ws5b0n0_53), .b(ws5b0n1_53));
adder_half ha132(.sum(ws6b0n0_54), .c_out(ws6b0n1_53), .a(ws5b0n0_54), .b(ws5b0n1_54));
adder_half ha133(.sum(ws6b0n0_55), .c_out(ws6b0n1_54), .a(ws5b0n0_55), .b(ws5b0n1_55));
adder_half ha134(.sum(ws6b0n0_56), .c_out(ws6b0n1_55), .a(ws5b0n0_56), .b(ws5b0n1_56));
assign ws6b0n0_57 = ws5b0n0_57;
assign ws6b0n0_58 = ws5b0n0_58;
assign ws6b0n0_59 = ws5b0n0_59;
assign ws6b0n0_60 = ws5b0n0_60;
assign ws6b0n0_61 = ws5b0n0_61;
assign ws6b0n0_62 = ws5b0n0_62;
assign ws6b0n0_63 = ws5b0n0_63;

adder_half ha135(.sum(ws7b0n0_1), .c_out(ws7b0n1_0), .a(ws6b0n0_1), .b(ws2b4n1_1));
adder_full fa876(.sum(ws7b0n0_2), .c_out(ws7b0n1_1), .a(ws6b0n0_2), .b(ws6b0n1_2), .c_in(ws2b4n1_2));
adder_full fa877(.sum(ws7b0n0_3), .c_out(ws7b0n1_2), .a(ws6b0n0_3), .b(ws6b0n1_3), .c_in(ws2b4n1_3));
adder_full fa878(.sum(ws7b0n0_4), .c_out(ws7b0n1_3), .a(ws6b0n0_4), .b(ws6b0n1_4), .c_in(ws2b4n1_4));
adder_full fa879(.sum(ws7b0n0_5), .c_out(ws7b0n1_4), .a(ws6b0n0_5), .b(ws6b0n1_5), .c_in(ws2b4n1_5));
adder_full fa880(.sum(ws7b0n0_6), .c_out(ws7b0n1_5), .a(ws6b0n0_6), .b(ws6b0n1_6), .c_in(ws2b4n1_6));
adder_full fa881(.sum(ws7b0n0_7), .c_out(ws7b0n1_6), .a(ws6b0n0_7), .b(ws6b0n1_7), .c_in(ws2b4n1_7));
adder_full fa882(.sum(ws7b0n0_8), .c_out(ws7b0n1_7), .a(ws6b0n0_8), .b(ws6b0n1_8), .c_in(ws2b4n1_8));
adder_full fa883(.sum(ws7b0n0_9), .c_out(ws7b0n1_8), .a(ws6b0n0_9), .b(ws6b0n1_9), .c_in(ws2b4n1_9));
adder_full fa884(.sum(ws7b0n0_10), .c_out(ws7b0n1_9), .a(ws6b0n0_10), .b(ws6b0n1_10), .c_in(ws2b4n1_10));
adder_full fa885(.sum(ws7b0n0_11), .c_out(ws7b0n1_10), .a(ws6b0n0_11), .b(ws6b0n1_11), .c_in(ws2b4n1_11));
adder_full fa886(.sum(ws7b0n0_12), .c_out(ws7b0n1_11), .a(ws6b0n0_12), .b(ws6b0n1_12), .c_in(ws2b4n1_12));
adder_full fa887(.sum(ws7b0n0_13), .c_out(ws7b0n1_12), .a(ws6b0n0_13), .b(ws6b0n1_13), .c_in(ws2b4n1_13));
adder_full fa888(.sum(ws7b0n0_14), .c_out(ws7b0n1_13), .a(ws6b0n0_14), .b(ws6b0n1_14), .c_in(ws2b4n1_14));
adder_full fa889(.sum(ws7b0n0_15), .c_out(ws7b0n1_14), .a(ws6b0n0_15), .b(ws6b0n1_15), .c_in(ws2b4n1_15));
adder_full fa890(.sum(ws7b0n0_16), .c_out(ws7b0n1_15), .a(ws6b0n0_16), .b(ws6b0n1_16), .c_in(ws2b4n1_16));
adder_full fa891(.sum(ws7b0n0_17), .c_out(ws7b0n1_16), .a(ws6b0n0_17), .b(ws6b0n1_17), .c_in(ws2b4n1_17));
adder_full fa892(.sum(ws7b0n0_18), .c_out(ws7b0n1_17), .a(ws6b0n0_18), .b(ws6b0n1_18), .c_in(ws2b4n1_18));
adder_full fa893(.sum(ws7b0n0_19), .c_out(ws7b0n1_18), .a(ws6b0n0_19), .b(ws6b0n1_19), .c_in(ws2b4n1_19));
adder_full fa894(.sum(ws7b0n0_20), .c_out(ws7b0n1_19), .a(ws6b0n0_20), .b(ws6b0n1_20), .c_in(ws2b4n1_20));
adder_full fa895(.sum(ws7b0n0_21), .c_out(ws7b0n1_20), .a(ws6b0n0_21), .b(ws6b0n1_21), .c_in(ws2b4n1_21));
adder_full fa896(.sum(ws7b0n0_22), .c_out(ws7b0n1_21), .a(ws6b0n0_22), .b(ws6b0n1_22), .c_in(ws2b4n1_22));
adder_full fa897(.sum(ws7b0n0_23), .c_out(ws7b0n1_22), .a(ws6b0n0_23), .b(ws6b0n1_23), .c_in(ws2b4n1_23));
adder_full fa898(.sum(ws7b0n0_24), .c_out(ws7b0n1_23), .a(ws6b0n0_24), .b(ws6b0n1_24), .c_in(ws2b4n1_24));
adder_full fa899(.sum(ws7b0n0_25), .c_out(ws7b0n1_24), .a(ws6b0n0_25), .b(ws6b0n1_25), .c_in(ws2b4n1_25));
adder_full fa900(.sum(ws7b0n0_26), .c_out(ws7b0n1_25), .a(ws6b0n0_26), .b(ws6b0n1_26), .c_in(ws2b4n1_26));
adder_full fa901(.sum(ws7b0n0_27), .c_out(ws7b0n1_26), .a(ws6b0n0_27), .b(ws6b0n1_27), .c_in(ws2b4n1_27));
adder_full fa902(.sum(ws7b0n0_28), .c_out(ws7b0n1_27), .a(ws6b0n0_28), .b(ws6b0n1_28), .c_in(ws2b4n1_28));
adder_full fa903(.sum(ws7b0n0_29), .c_out(ws7b0n1_28), .a(ws6b0n0_29), .b(ws6b0n1_29), .c_in(ws2b4n1_29));
adder_full fa904(.sum(ws7b0n0_30), .c_out(ws7b0n1_29), .a(ws6b0n0_30), .b(ws6b0n1_30), .c_in(ws2b4n1_30));
adder_full fa905(.sum(ws7b0n0_31), .c_out(ws7b0n1_30), .a(ws6b0n0_31), .b(ws6b0n1_31), .c_in(ws2b4n1_31));
adder_full fa906(.sum(ws7b0n0_32), .c_out(ws7b0n1_31), .a(ws6b0n0_32), .b(ws6b0n1_32), .c_in(ws2b4n1_32));
adder_half ha136(.sum(ws7b0n0_33), .c_out(ws7b0n1_32), .a(ws6b0n0_33), .b(ws6b0n1_33));
adder_half ha137(.sum(ws7b0n0_34), .c_out(ws7b0n1_33), .a(ws6b0n0_34), .b(ws6b0n1_34));
adder_half ha138(.sum(ws7b0n0_35), .c_out(ws7b0n1_34), .a(ws6b0n0_35), .b(ws6b0n1_35));
adder_half ha139(.sum(ws7b0n0_36), .c_out(ws7b0n1_35), .a(ws6b0n0_36), .b(ws6b0n1_36));
adder_half ha140(.sum(ws7b0n0_37), .c_out(ws7b0n1_36), .a(ws6b0n0_37), .b(ws6b0n1_37));
adder_half ha141(.sum(ws7b0n0_38), .c_out(ws7b0n1_37), .a(ws6b0n0_38), .b(ws6b0n1_38));
adder_half ha142(.sum(ws7b0n0_39), .c_out(ws7b0n1_38), .a(ws6b0n0_39), .b(ws6b0n1_39));
adder_half ha143(.sum(ws7b0n0_40), .c_out(ws7b0n1_39), .a(ws6b0n0_40), .b(ws6b0n1_40));
adder_half ha144(.sum(ws7b0n0_41), .c_out(ws7b0n1_40), .a(ws6b0n0_41), .b(ws6b0n1_41));
adder_half ha145(.sum(ws7b0n0_42), .c_out(ws7b0n1_41), .a(ws6b0n0_42), .b(ws6b0n1_42));
adder_half ha146(.sum(ws7b0n0_43), .c_out(ws7b0n1_42), .a(ws6b0n0_43), .b(ws6b0n1_43));
adder_half ha147(.sum(ws7b0n0_44), .c_out(ws7b0n1_43), .a(ws6b0n0_44), .b(ws6b0n1_44));
adder_half ha148(.sum(ws7b0n0_45), .c_out(ws7b0n1_44), .a(ws6b0n0_45), .b(ws6b0n1_45));
adder_half ha149(.sum(ws7b0n0_46), .c_out(ws7b0n1_45), .a(ws6b0n0_46), .b(ws6b0n1_46));
adder_half ha150(.sum(ws7b0n0_47), .c_out(ws7b0n1_46), .a(ws6b0n0_47), .b(ws6b0n1_47));
adder_half ha151(.sum(ws7b0n0_48), .c_out(ws7b0n1_47), .a(ws6b0n0_48), .b(ws6b0n1_48));
adder_half ha152(.sum(ws7b0n0_49), .c_out(ws7b0n1_48), .a(ws6b0n0_49), .b(ws6b0n1_49));
adder_half ha153(.sum(ws7b0n0_50), .c_out(ws7b0n1_49), .a(ws6b0n0_50), .b(ws6b0n1_50));
adder_half ha154(.sum(ws7b0n0_51), .c_out(ws7b0n1_50), .a(ws6b0n0_51), .b(ws6b0n1_51));
adder_half ha155(.sum(ws7b0n0_52), .c_out(ws7b0n1_51), .a(ws6b0n0_52), .b(ws6b0n1_52));
adder_half ha156(.sum(ws7b0n0_53), .c_out(ws7b0n1_52), .a(ws6b0n0_53), .b(ws6b0n1_53));
adder_half ha157(.sum(ws7b0n0_54), .c_out(ws7b0n1_53), .a(ws6b0n0_54), .b(ws6b0n1_54));
adder_half ha158(.sum(ws7b0n0_55), .c_out(ws7b0n1_54), .a(ws6b0n0_55), .b(ws6b0n1_55));
assign ws7b0n0_56 = ws6b0n0_56;
assign ws7b0n0_57 = ws6b0n0_57;
assign ws7b0n0_58 = ws6b0n0_58;
assign ws7b0n0_59 = ws6b0n0_59;
assign ws7b0n0_60 = ws6b0n0_60;
assign ws7b0n0_61 = ws6b0n0_61;
assign ws7b0n0_62 = ws6b0n0_62;
assign ws7b0n0_63 = ws6b0n0_63;

assign out1[63] = 1'b1;
assign out1[62] = ws7b0n0_1;
assign out1[61] = ws7b0n0_2;
assign out1[60] = ws7b0n0_3;
assign out1[59] = ws7b0n0_4;
assign out1[58] = ws7b0n0_5;
assign out1[57] = ws7b0n0_6;
assign out1[56] = ws7b0n0_7;
assign out1[55] = ws7b0n0_8;
assign out1[54] = ws7b0n0_9;
assign out1[53] = ws7b0n0_10;
assign out1[52] = ws7b0n0_11;
assign out1[51] = ws7b0n0_12;
assign out1[50] = ws7b0n0_13;
assign out1[49] = ws7b0n0_14;
assign out1[48] = ws7b0n0_15;
assign out1[47] = ws7b0n0_16;
assign out1[46] = ws7b0n0_17;
assign out1[45] = ws7b0n0_18;
assign out1[44] = ws7b0n0_19;
assign out1[43] = ws7b0n0_20;
assign out1[42] = ws7b0n0_21;
assign out1[41] = ws7b0n0_22;
assign out1[40] = ws7b0n0_23;
assign out1[39] = ws7b0n0_24;
assign out1[38] = ws7b0n0_25;
assign out1[37] = ws7b0n0_26;
assign out1[36] = ws7b0n0_27;
assign out1[35] = ws7b0n0_28;
assign out1[34] = ws7b0n0_29;
assign out1[33] = ws7b0n0_30;
assign out1[32] = ws7b0n0_31;
assign out1[31] = ws7b0n0_32;
//assign out1[31] = 1'b1;
assign out1[30] = ws7b0n0_33;
assign out1[29] = ws7b0n0_34;
assign out1[28] = ws7b0n0_35;
assign out1[27] = ws7b0n0_36;
assign out1[26] = ws7b0n0_37;
assign out1[25] = ws7b0n0_38;
assign out1[24] = ws7b0n0_39;
assign out1[23] = ws7b0n0_40;
assign out1[22] = ws7b0n0_41;
assign out1[21] = ws7b0n0_42;
assign out1[20] = ws7b0n0_43;
assign out1[19] = ws7b0n0_44;
assign out1[18] = ws7b0n0_45;
assign out1[17] = ws7b0n0_46;
assign out1[16] = ws7b0n0_47;
assign out1[15] = ws7b0n0_48;
assign out1[14] = ws7b0n0_49;
assign out1[13] = ws7b0n0_50;
assign out1[12] = ws7b0n0_51;
assign out1[11] = ws7b0n0_52;
assign out1[10] = ws7b0n0_53;
assign out1[9] = ws7b0n0_54;
assign out1[8] = ws7b0n0_55;
assign out1[7] = ws7b0n0_56;
assign out1[6] = ws7b0n0_57;
assign out1[5] = ws7b0n0_58;
assign out1[4] = ws7b0n0_59;
assign out1[3] = ws7b0n0_60;
assign out1[2] = ws7b0n0_61;
assign out1[1] = ws7b0n0_62;
assign out1[0] = ws7b0n0_63;

assign out2[63] = ws7b0n1_0;
assign out2[62] = ws7b0n1_1;
assign out2[61] = ws7b0n1_2;
assign out2[60] = ws7b0n1_3;
assign out2[59] = ws7b0n1_4;
assign out2[58] = ws7b0n1_5;
assign out2[57] = ws7b0n1_6;
assign out2[56] = ws7b0n1_7;
assign out2[55] = ws7b0n1_8;
assign out2[54] = ws7b0n1_9;
assign out2[53] = ws7b0n1_10;
assign out2[52] = ws7b0n1_11;
assign out2[51] = ws7b0n1_12;
assign out2[50] = ws7b0n1_13;
assign out2[49] = ws7b0n1_14;
assign out2[48] = ws7b0n1_15;
assign out2[47] = ws7b0n1_16;
assign out2[46] = ws7b0n1_17;
assign out2[45] = ws7b0n1_18;
assign out2[44] = ws7b0n1_19;
assign out2[43] = ws7b0n1_20;
assign out2[42] = ws7b0n1_21;
assign out2[41] = ws7b0n1_22;
assign out2[40] = ws7b0n1_23;
assign out2[39] = ws7b0n1_24;
assign out2[38] = ws7b0n1_25;
assign out2[37] = ws7b0n1_26;
assign out2[36] = ws7b0n1_27;
assign out2[35] = ws7b0n1_28;
assign out2[34] = ws7b0n1_29;
assign out2[33] = ws7b0n1_30;
assign out2[32] = ws7b0n1_31;
assign out2[31] = ws7b0n1_32;
//assign out2[31] = ws7b0n1_0;
assign out2[30] = ws7b0n1_33;
assign out2[29] = ws7b0n1_34;
assign out2[28] = ws7b0n1_35;
assign out2[27] = ws7b0n1_36;
assign out2[26] = ws7b0n1_37;
assign out2[25] = ws7b0n1_38;
assign out2[24] = ws7b0n1_39;
assign out2[23] = ws7b0n1_40;
assign out2[22] = ws7b0n1_41;
assign out2[21] = ws7b0n1_42;
assign out2[20] = ws7b0n1_43;
assign out2[19] = ws7b0n1_44;
assign out2[18] = ws7b0n1_45;
assign out2[17] = ws7b0n1_46;
assign out2[16] = ws7b0n1_47;
assign out2[15] = ws7b0n1_48;
assign out2[14] = ws7b0n1_49;
assign out2[13] = ws7b0n1_50;
assign out2[12] = ws7b0n1_51;
assign out2[11] = ws7b0n1_52;
assign out2[10] = ws7b0n1_53;
assign out2[9] = ws7b0n1_54;
assign out2[8] = 1'b0;
assign out2[7] = 1'b0;
assign out2[6] = 1'b0;
assign out2[5] = 1'b0;
assign out2[4] = 1'b0;
assign out2[3] = 1'b0;
assign out2[2] = 1'b0;
assign out2[1] = 1'b0;
assign out2[0] = 1'b0;

wire low_c_out;
z_adder_select_4x8 my_adder(.a(out1[31:0]), .b(out2[31:0]), .c_in(1'b0), .c_out(low_c_out), .sum(result));

wire [31:0] up_sum_0, up_sum_1, up_sum;
z_adder_select_4x8 my_adder1(.a(out1[63:32]), .b(out2[63:32]), .c_in(1'b0), .c_out(), .sum(up_sum_0));
z_adder_select_4x8 my_adder2(.a(out1[63:32]), .b(out2[63:32]), .c_in(1'b1), .c_out(), .sum(up_sum_1));

assign up_sum = low_c_out ? up_sum_1 : up_sum_0;

wire [31:0] xors;
	genvar i;
	generate
		for (i=0; i<32; i=i+1) begin: loop2
			xor my_xor(xors[i], up_sum[i], result[31]);
		end
	endgenerate
	
	wire [7:0] xor2;
	generate
		for (i=0; i<8; i=i+1) begin: loop3
			or my_or(xor2[i], xors[i*4], xors[i*4+1], xors[i*4+2], xors[i*4+3]);
		end
	endgenerate
	or neq_or(data_exception, xor2[0], xor2[1], xor2[2], xor2[3], xor2[4], xor2[5], xor2[6], xor2[7]);


endmodule